��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�F����c8�@S�B�v�Y��`E�.�}j'.��ʠN�r-���fϔa��/I)���'����-&3��"�SO�5��J�V;A9..M���Z�ΨW<r��v��\AZ��kO����ٯ[n���g"�2t�����1���v`iK�M��j�������_��&�Ҹ ��S�)=MB�k݊OH��n��]��/ge��<��Om2�"ˏv�`��ľ�"Vϼ�����F� 6� <b�%�It�b���E@q+��ۦ��bڇ�ߙ�i�������{eq
톟�u�#�*��ܰ���ev!M&�)4J�ug�����ߗƺ# ���9B]�ȖWq�ڙ��a�m�������=MX�4�桹k��f��*t8"s��S�Jĭ�g�g���A�B��O�"��+�f��7e��d��͍깊v�ϤP�1��:��fi(@���O�]5���X�͎���� :��d�'\A��^S�] �d����T�}w��C�(��2�q��BB�z�n.�Rj|�Im%����R����(�+1	��(Bd����Q�����PQYl��<�ʅĐPKo#W��h��ַw��`�	t�o�G��( ����>�D����[��3��\L�/^����A ȃ��_Oe��>�t�t4��[���L_b *�r���8gb���g��� ���o��T�Π�7���#&�ײlC�}�"؟�9�z�����WҺN�*������"XQ�@/x�x��6���Rc�
.�Kx����΢h�;��YL�t��f녂�*����?��<�.f�gsS���NB6����e���U*k�w�&G���U��xqw{���ӎ���32;Gx���:��B�.9�B�nJ���9?�ߔ#&�O����Zjd��d�Wz߅�OlKG�������^y_�?o���&p)Z<H�Oj1u��p:�=��^�!����>�.�P�	����)�A�ɲ�ʵnf��ss���\5��h����7`O��[�u�j�v��uv�,�O�����Ϗ�7��`L�8�)���d���Ϥ��+����S=}��q�J�WRğ�\;_զ2��Q��D��*���x��5�[ޏ?V�J�w=(����O}�JV�	�a9�B`׼��4�j([�p.9
l�r]�^E���B�}��n�E��|ᥕː�$���"=S�	�]+���Ifny�b,>�s��<Cf즻?��eY��R�`�9��.}�{������f���KO����q[�av�g[�V;�E�Y_:?��z�\:]�Jض,�w�`�C��s�ld� `��i�h�|F�<����N7 1�,�g��5�)�8U�qhL�Z������9\w��R����e��}q�����.3S��w{!զ�����
� �Ā�t�s����.U�� 諟�x�t�F1��҃uQ�%;	lӰV�ڛ��o�s
Rz]9K�*�r� ����ʞ����yr���
ۋ� ��]t�mS���#b7�|�J�XSu��A��2��Mcen��{һ�$,��s&Ë�t/�[&�pط��&�R*����3Wx�5��uMXW�&*K�	A�P�����9����k'--����	k֚�q�H��	<�Ӝ`�.;D�D��cc�4�H�:r�{��í���Fc�)8����Z����Od���Q:��Q ^�+�P�z*/-~�����m���ղ�
S���� ������HV���O'��׸v�91�K�����R���m�H�]0�d���2�����EMB^� Fbb 94���q�(qb�sTq�k��f��

���j�YE�?��h�S���.^�:>"�Yv���Z�^�d'�FW��
2ʒ�L�J^@A.�Z�Է��y� 4�T�^������=ﶳ�����5QO�&�:t~q/B-1+zz	���5��-PK�G�ꈗ�@��CiL�S�#{Ԕ���y�Q��o���p��
�) ��>&��z�g#T�(PH�'\�
���x�j
�����ޤ<����ӲD����R,��~�Ѓ����!`&�#`���ߤ�_3�N��E6�o-�Na�>xCN۝��,����	2xQ������Ms�E�XB�Ć�* �p)�Q���BWW��,K0�tK椴$��bK﷋�X7�=WKI�ObZ���W3`g�"+�m��?��Ij����ܥ���B�$M�O{qf8,\���br2.L������>�~�aj�v�o4���n��8^��oDq�І�r�8�O�Զ�g*��/�;E>�����rn�Y�@�/wrV5�sv��4�L/�h ��X��Q���n��0N)�Et� [��x�[Wr��m�aȑ^#/��B�5/C;���a�9Q�&�kFH9�1wh2OQw2fz^�� s7���k[�(��+���+��_����qX�6A&y��c �&��;7�;Jޏ�:)�@�\K ��F�R��9XB���k����W�������-9ʔ~���[qp=5{T�:��&.C&��d����@�j�}U�u��?�bW�B���LUPq�O���6?��?�r��O�����h�*j��Ʊ0�IJRw��� ɸ@�暐\sv��L�G`22���{����h�+��b���qg짦@�z�S�"��Iu�"��Gs�wY�ToH�;�� g�Ky��B!y��-��&6*ə��Ǩ�*����QÕ�t������Ur4�=�# g޹J֪�T�%U�)��<`T^s�V �Dq�H�iWb�{���A[�/09���d�ӣ��ER!�R��a�XQWu�TMҫJ@H���o������:6�~'�1^�ʨ�-D�1Z��B����r��x�!����7�6��2��VF�� ��ߑ�u�Y_�����lZ�\�|�F��;�/�%%+ߵqt�(h�tɓ��;�S}9psmc2����W�Rvһ��P	i���W!�N�(�M})C��6�ۂȾ���.�˅I�~��<~��J8�l����8p~�w.w�r��^Wo��'Nޡ^��HV�1=�쿤X�Y��lDL�E���}�IhQR�,dQ�@�#$�򫠻��}%�h�Kۃ�S�TEy�	�U_�n���{#-"� I^`K�}��9P�1+.VBHe�N��r~~����aA����w����N*���&���/h�$ټH͘����H��|d�e|2+&��qeu���B�Λea!#'3�o����=3�����(����x��	[�G�ě6 �B�W��fY>u�Kb���b�Ը�LQ��X�u������#&-�yo��{mIUkZ&��ʆ~�k�0���qc��)���c!�c��b�m�H�[}f�Ќ��Nҩb7���O�d��� �@c/�5A�CQZHa\��u`��;c	�̗���D��8��m���^ő��N30Qs��%f��2��˾�=�2:��i07����WϤ\�%�����O�kUC�%kd��0,���ߑ�=�./9����V�׻��{�5��h�,'蹋S|�ŵ��Fcf�p���F�������=�#�D0��V��Ƃ�Q����{[h<���S��)X�"WZodM�G��&v�fs�]t�Q���`~�GC<Է<���1[���g �|g����Bۃ��X��H~w�,���G�F�?��{	�[|�O2���6�|���*���2�R�c�c�L�AB�w]�� �|��8�9%�)6�xêM��F��P��Տv{���2 "������%F���yM+*��T���P�0T�؆�9�������Ǽu���R􆡨Ƥ�x�a1y�xN�`˶�B�~��%	Y��;B�{߉V�,g�9+;[AЄ7�$G�^��*#�-)g�{�9�K�S�X#�~e֐8���(v���H�}�u�ǈ`��Ci�ܖ�	9����8�z>�p��s���I�3ZlLv�l�lS�@˄���xeL����jF���`���(����b�6QU���)�K� [��H�i��E-��]�N�^�R|H��s�k[�mO�'c��#r���^٤C��8��p(Y�i�m�	�'�w$^�QB&�y\� xķq��M*���7+y�q\����,lܝ9�����g�l�.����|���<�:v<	΋7�̂ܥ�C�"-K0 �^g3��;/���4":C��?)2|Gg�%C�� QE �+<��'�����O���y��w�z������*OE��ቤ��U�1 ��}%����;+�3�>���"�C���}�u��mϊeTT�pv�}X�*?���T���v9����zb�Fa���?��h�����S$�e�㦖�� �M�48�.�u��;[�V�ԝ	������$H�P7���`t�q��^��] �׳�I�7s�T��K^��}4�NA÷d�J�#@�K��a�u��-��1N�g�ݻ���-�zx�{c��1��|D�*K�h����夼�5='�H�tDĉE<~�˻�>�l"ʢ�_g��v�0���sF�P{߬6�y<��9�fk��!���;��`��F{�3
k�B�gB����R�C60Ǻ�0��E,x��)����f��̼�%x^�=�(L��FX��dQ4��'/Np�4"�E�z���,��ۘcZ�����3h��
�e��p�H�x���P��3Ĭ����_|�K��8z�M�g�;�)��A�DMs}:�>�u�Uޤ����u�ǁ�#�m�q� ���<�V�(��&�������rC5,���P��ݷ�Pc���FE�ly�w��f�3tfZ�[ae�G�̫=����e�>� -�S�=�M��!�#�X$��H�H�#0;Q��w�ef��#V�s�Ngc��H�
.��Ly��[{������e!8��w:��e�з�4��cz��~� lK��a���Z"�qy�Ȱ���B9HU��YDB��B���:.���)Y =�i=�[b��m�>lo`�' �n�I"���dS����[�Ύ��4%f_�W{WO�D~4�'�:�އ'񋄣���d��l39+��;Ȣ�}�T�UCi��Q98Au��"�G�YT�_w<���j�g;������F��>�QW�J���5O��g�,��B��=��`O�L|?�5�csXvVs��I����V�/�p�tc.��`t��bh����m��|�J�
+�e�Y�ĩ�2�piV%�r|G9*�k�	��?�;G��9�K�T+�R8�I4��kƎt�33b��8w��9�ϒy'̍��[vg:L�RZj;�($�7￫�~ɡ���TC+k������H��g����1 !w�Y&�Qғ7lk�pi�G��C�Xc}3��;�"L `1*��o�M��0�Y����Ӷ��W� 7,��w���0!��{߉A�Z����!rZ�d�DP�0��� J����P	%h��$�k�L;"�'d{qƫ��vu9����	��^3�tibqEX�ܮ3��}������)�ŭ�/42��z��5�u��|p�Vl=\�@�I��;�B�AٍB�7�	�N#=��Y��y�� R����x`����� 8��cjƝk؄�E�wk�'��J����|
N(��8 �����u�uɞ��� �� ��pI�xր^ъ
����D�8)��SX=E��$ ��!T�����ѝ[�3�Xo�Y�Y�у92����,L��5���"�BGn�{���YrS�j'���R���xk�xh��I����j~sIwE,w1ƫ�=6g�Ԕ���p��,�G`�U�/��咥4�r�~�Z��	��9����"Q^�^=��C�aXHI궸�L}y�/�^����c#�#���YCv��γVȫ�-O@���
Nwv=:�h�,�*�5�������ƹ:3�s5�:mC�Z��*��"���'!n�šp�s��4�a�{.��h{c
��g-��A�̇H���*"l�][��33M-8�
���%�(C��J?f�A2_桓m�-�=U�m�����S�\߀o3�ʤW�9X��x ��(H��Y�����$�[�B���� DC�Ea�a�tu=h���s��0��NE��x��Rb0�׶�j��jyp��9UY��cI����z�q��n%��@#4�}V7�*�dX��a�c"A<B�9���R�&�Vs#���#�D��k^?l��5�06K��cc�<$B	�1��+��'
ڥ�rPS�V�7����B/K�Ww����\����"�
����J�Mud��o�� 5�����H	gJ=�^�# ��ه��^M)�5���vP����h(��oM���
sI>Z����lW��jD�h���u8D���\�l+*H��=½�圭',��� �� ޝ>|ptpj�U~��`�5hl5"��ϵt+���y[�oX(L��\��b�����k�/1*J4^	ey1�g�32b�!�4���<l��{Ĵq�p	�^�9*�L��8	��ΣA�L#�HoCu��j!�7f���B\�$>_�ߡ�a���!��^>W���_�z�"
��,1;)ma