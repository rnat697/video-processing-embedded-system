��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P��A�?��cܑw��=f�������fl5;�7�q��Cªx���K��O���y�Ȟ#�∁.��r��;D��N|4�ʔ��-��ܖ��2��iʕ��[������eF.��'f���B�5�=&��fTa3^VL�[�n��b �g���u.`u�zZ�'9�`��,�y�]x�3|����һ�{�>��)Sӫ\���AeEʹg�DF��SF�e�~�2�����MMyn�k�Dw��wE8H�D�DfH)��W��ZU����Y�{J�v��G���t���z���O%��������s�I�:�?�z�#wƦ�:oX����*^\(�X�j�S �ē:l�Pa$�|����28�P{P��6�3���T�$ـTG��{��T-CR�3�y,�R�;��R��Ǭ��Y�G�J�ר�Wf�2��;�ܼ���7 ���%Zm��;�����O'�JV�[1��4-�O�j@J{7ג�MA����^���:��IB W��������A�t휁6����$� 0�Jb^���2��隗Tk��Ϋm�&��2rU�q��( �����]�3A̚iEivV���>�F0���9AO�C#�[?��og�fyp�r0gV���E��(&�S����$�9��ypt;��(��l�L�c3/]�r��1�����U�ǿ��
R����T(�:�W6���*�� �Zlu��T�����=���ȿM]�� �S��;�[� ߼�f�X��&�L�^��OB'�]�؎[f�$�a(�����ad&�c!�**s��͚t�km�b:x�$-���۳�`��6����z�H�Aǧ2#NY�N9W��Z��,�q}��l��yR�����P�

l��[~R���Q{�1�&#~lܱ���b�l��n���	x#���m��=-�v���݅\O�(�d��J�zI�t����z���űaj-���X�K����8dv����h����V1����4��>(�K��� %��&6=�`(<�/zrK`R�:�0b;x�&A����jF���q dr�!y��=�5.ـ�j��.�P��������u�]���V�V����!Rx��x�	1j��Ŧ8BQ���9�wZ�/b�ۙS��]�*�JWD�܋F�r����ۧ�i�r�f*�j��Fuj�]�?y}������e�X���xF"i�4
_-���j	�[�1
��9�cO��[�Y[en���@G�#_?�c{��4�5��e���}2�E+��P�]��(�m���5׎�4��;aO���o�ؔb���c��H&Ϲ1֡�#3P��qk�ꀡ�H,ҷ���q�+��&��-`�ѱL@��!�!n�2���+�n���X؁�H���"N#���o}�0��0
N ���r���Z<�ڥ�ұq g����"�bAk�Z��b�\j��?`-�)�������Ļ;,)(Z�k�2��t�����R��:�O�e�W���,�a����D�{�����MYr��O����{nF�"�#PT���Q��<л���&��'T����*��w0��+El�i-�s���z"`ɻ��S.�s��x<�H��Z�lQY\QGkWm%b��#�����=,8��L���Fe�n�3"V%
��,���h��-P��&"��qJn����~�S]ތP��N���`����i����DnF�@^�f�IN6N$w����?��/���ı��D��D%V	�@����(�y��8��!Aui,
]�0g�Lm���_So����k�AI2� j�qhڿVN�-G�D'&�mI����8�8�B�4s�+�;����`�jjqc>]Z�i� ��.�f9n�A?M�c��-:�Z\�;��%��Ҍ�7w���5�
����vH�d�؆?6���'#;�l�;���s1JVfDwop"<Y��'�ǃ�>,
9d�E�@ߴ+_&������kV�����%'g�T��F��s��G����y�;�K�Z]�,�&��n+\sc�'Q��{�51�cݨ��%��N���ZDC�Y����lыʹ�K��޹5Iֵ��#2F�JPCVA�&qh\����.�Y�;�?�����E�>��WZ�� $����5@xg'����Bjy`=$ٺ	�	h6C#��1~�ۍ㚍%�\.����+�$/?r�-%w����f��۪\>D�!��J���Ĺ�_�
q5�5V����'!p���X�X�㠅�?�����փz*͋����}��+jӚD�������A)��o�pF=�N 
��n���=ݢ�{~��5�A�Ë�4��O�-�y����Gli�-J`�{;����%k����oz�����\��Ke�\�+��� 9��>�sю$��A	Liݵ�BD�J^����O>
�]w؉���m.�S��T>��<E�(;B���ܼ��:8��L�?O� �Hbhd�Z|XFW�1to����\2���纗kq����щ���9s�v��ݨ�xʢm�"f'���K����#��w� �!�g�sqNK$���뾄�$P]��8P��d�N�*���N�o�0.��v�t���39Lt�����M߫��jT�[�| I����\�'��D��j�O�M%��yu iw������/D�3��� ��ߒW�1P����H��#�~�z���o �|^�Ě�F|�F���V�z��,!Q��5���l	,�-�v�|6��=B'��z@O,Q��z�T���X.u�G6{�~����({�va}��&��/9(�z�Mׅ����:�vM��҂��#"%��R�-J��y��7�֨Q���>�pv���m�l�ě�]]�g��.FO�ŷ�N��cO&�\@"�QH��@�u+����)�P�&���q��<����%���-F���HZ����u|,�(OI+��ױ'F�,�+��`q�7=�2�����a��5B�,�g��/�[-�ҨB�����SP�M��H�*|�)0�*�l�y~�=�L�&�zűG8�a���{��;�g�e���4rBR�`�-���M�U,���yI��}s��a�T
HNv��9n;A8�ȿHD��H��A�_Ku��H��gX�Q�Z�ʥ��v;jJ^(�}�aVC��٧-��_̯����4���G��c�2�8�n�t�X�T�,`!�]����'=\��)����+���C�QR'fy�շ�c���:j��D� �6[��BM�Q��M>z1^e
7���؆� k�8y���9+�R���.�߯�J��}�a�zzV��k���Dҭ��%����,ڦo�dI�-���5��{V�4�>=�����@&��6z��-�u�,ې�� �!��0�9�fKɸw=}�G�Ą0Y\d(u��f���ˑzl��Җg�j��"��Sn���m�/��s;D\7ifY/|VU� nI��_�.�ќf��#���c��rz�Y�䜸 ��y0�, "ђ�Ef�M������w�]�)���&����A<�6|o3D��i�s�f��Ⱥ����XW��][�>��!T,7�DN�Q�������&6���?=Ƃ��7�A�5D��qe��eR��}O��Ok�E8D6�۫��&g��֢�p\���#o���I��[hSc���sȚ�E�o���W�7+�=���RE��pk]��%���$nDخ�,���xyk�
x�^#��|��)��)��"���!��k��)��T$�^�ܲ���E�o��n*]��c^��E�}	�O�)��F��Ț���L����f���q���#_���%f5�4�3W�+h���a��rOo!J4�I�ؽ*��"�g�����Ȋɹv���Y�q���c�/���Z6;�r���&+�fߩ��������:�i��Vʷd�$ ����w!5��9g�k�y(�<��&A�N�!��H�o�?��ŧ%�$�|��([�P�_B��	����nm��ϔ=��b�eѯ��m�?�*��k>�z�O���� !��%K��-�p�\DwR%}�$͓�I?���~�Ͼ�ph�b��1H9������	qڃ U��S;��G"L���Y2�[�����Q��p����w(��~��=F*10g.J���r�p�ӽ���5�`Y�Zz?Z��-c#8o$��A���s1�
�a�Z�U�"v������aN�1:��m4�ê�|π��Q΃ʑ|��,/];�h�eG2�@d��?�J�e1�#n�S�8�]���o��2iZ%���0]����N^+���r/�:��X�k��[<���z��LH�ɺ��6o���H&/-<�G��/5� ��npvM�%�{�m\(��cP�!��g�ŧ9�&X�G��U�*$��=��W�8�BA
��3�e���.j}f'�M����"�iO��R�cB��[��0��˝��̦�ڗp~�	�dL֊�F�_��;2�Ԝ��~��˨Ǔ��n��7����Q~���p�j�+�W��Gx��g�u-=�2��zэ���"?��fْl�H7��g"op��(��=w�B�X����z��O�'�Z�S��""EP�/cx���Y�N�e���dK�MA��*�M���2���=u���D���Fz�%��4��R㤪��w�Xs�<]�h��ߒ7�i�7��YܷeJ�)�FО�4�:|?{1$qܰ�d�-���Y���+��M�݈>�ų�ch"���h�3^P\~��+Y����~]$�����J:R���o�Im9#�X�ϓ�:��Ҁ�KQ�,����H�p�*%�Nǈ�r���Z�Px7����6�
�IK8�^:�w~�O����IG��4~��(ё`S���R�`��/�S�kf)��<f��t�
>��Ugy��1�<r�V�^��yy�!Ú�ֹ`h丒�[�}ݓ��حД�B�����d}�P�Xє�}��x.W�t�s��p����5SU9V4c2o�$�*�Z~�.F�J�%��,��m�R�!�-�Jm���V��ұ�Ct�G�g����b8���`M^y0U���G��tc�C�%H
�k����<b�^��{��ɇ��=������|	���<���Ӝ
�OV�PUW��%�if�i�cmO�_���4���$K)OO����z�r��`�l? ���~�[����X6`g��l�4�wΥ
�"�M��InWK�yef5Vs��Đ\��|�ֿ�3�>y4�|&��m�j8�*����O�*ݺ��=��-�C�eQ
��W�+�s��9�h�s��R�x7��\��A^��[�O-���Nu�8�����
�3�:ғ�7I�\I��19����L�c��gt�(�W}�j�,��!
Ճ������t2�����^�6��5R
���z����a�$%�"�,�^�z��2�J0��X���:�|mnSX�ً,�۫p�| ͆���}R�ˋ�|�d%�>9���}m�~���wJ� ��	��%�G��d�붫K�SL��HN'�0�k���5	��Tg��
@��nG�~D$��&��ʇ�o4�c��!�bٽQ��\4r�o�����Z׭�2���f@����3J��ʠw~W���7E��66C^�rqbVU�����:�Y������)���|@?��� ��5[&��O�W?���:J���Gg�����ӐF�/��-�q�+y]p��3��_X���R��k�lE ��7{EN�j�7q���K���	E6�Ch�&(�������~�kJ�{m��}�o��/j�p���Hxe�o�.��Xa���nܴqE�o0�`�c��K��Q�l���Q���%����+g���S��7���-���=��t�$^�yLaQAJ5��.^e�T�8��-j'�H<�Q����f�k>	�u&�aY�Mf��dU����B��;�0ZV�v��ֵܰg`�z�k�R"�Zm�$�RXٿ�1m�Z)�V�fܕ1�6�T�qu ��FQ���?뿡D[4�;�喘��Z��owk�[ L!�H%1<���{��S��H�(=O�����<��Q3�A�c���m����ڬ2����Pa��yv��L"��4��=�x�y���7��>���u'T+�Tq�F�kZ�N<��33+ͣ�AT����Am!�r(\p_��§��z ]�d�1(�ƒ�=��.h�p]U�*
����^��V�.�t�.6�T�h{��a8�I� 
���WW٘�J�<Ѱ�sj�u�%n���("�I�5�Mw�_Ox�~�V9���3�՗��_�v�,U�?S�}D�]�l]�W2	��^���zw��{k:���酞`d���oYjդ�4f܃�3�^@��ܲd0�����ZN��9�͍������~��:+E���zp�����\���z���b�-���H[)
A�VѭO�oL�f�
b�1��&C��n6�&�c���������so�Q|ܓ��i���M�Qa<���0�:{+B�7�:L���#�r��x�&7rW�4�qݷ0�����E��A[��%��b��q d�46B�q���>�Wu���u�gcf���o{A�!�V�j��3�L*5�킚�]�9�#�D���/�t>H�K�ф�ˊs������I[�j����Zy ����+�(��::�BKP#��.z�2�w�!j�b5怩&VC�F���(|���:�Bl`�����ݘ+~�W^@?�A�&�9_N����\C�6Ї���z0��,h������1K�c].���c���<>��Ij'�;�v0��{�CU��"�,�"���e��#��KBR`��2'�NF�̢v��	���&AZ�zƍ0_��t����bʶ��;3T� g"4Sp�}A�39A�-�]�r���$Wܛ_3:�vEs�Z{'2w����u��8���M�q=���ĉd&�q��|��ЦMc�#�c-�|^=jU�g���1�k�鱭5� 1����mM�s��{����.]�� �o�w�Wϗc�*9"�=���h������8Q��R�O�k�����T��)=���2c�[㦥?��?�g�����J��tȨ�,�����1_@+ٜ����O�=q1+T��5��z'��I�^�����5V]Y쳳��86;r(fq���6ӎ��=D��p����}�m���xJ�g�s��A����s`r��iX�	�D;.�;�xj����;,��ĖT�nђ&�gu�CѬ4���p�1�]ȫJ2=�\��\7
�HY��$Z�BY�#��@t%$�#�T pVTZ0��lZY/&���y|]^�d>Is�ƹsoI�.����R��e�X��iA��6fWb8."|&^���O=�)��ƙ��:�d�2�%�L�]5o��Hz�hd����� Gf�c��Pn��~=�NM�ޑ�G���?�[�H�TW�w���B���+y:�d��]�4 ��H՗p���ȃi���6QT#y�Ώ$Y&�[cI��5��[��i��:I5m	�ė�SjZ��|�J��ޠ�)���I��YH��Q7���/�a�X����6�}QS��_�g��|L3G��?�mF8�����A�;�tA�� ��P�q�F>/4�%Hl��83+ں����.V|�C�XɁK�p}���6�sć�@gD�)��A��X���'�]G(��\g��r�a��Ӧ����g�w`��5dٰ$�:]�cE0#�䞼LH�A��Ԫ��-?{���½��[�����mP@�t����^�k�摇O��T�v	^ɵ�R̯��X9��G)�����(>��׳���ތ�+��} ?B�+��U�@�AS ���?�ݲ�����b/aF�b��߫��I }n��v �N����9�+��wЕ� �=�G�Λ�$�	}M���s��q�bs0���`7 �`�]���m�,07Z�{;����b�A�KA��P\d}��
k�ls��g��@��O��djm��T[�1�L��)�pء3ڑ7Ez�gc�(��Z��(!��	_��=^�
�WF3m��d!g����*��bs�H>������ER�¥��>��ϩ5T)������4s��[���XfxH@<���6mjq������L��ԝ-�r�,�k���,��:]�jx,���f���2'?1Km#Ƹck!Dû����|����7�7���FS��4;�� ����'�����$a�pw����{����ni�m�c�5gG�<�X|	�m�!�mد�G�AV�)W,TW�j% ~7ʋ�'��9o�ϳ��S9��h��q:�� ��I��m���O�z�Pe�*�s���"r��C�t��<��ΊTe��CLt�2��J&�SI�6���D�:�+>�)�^d
�ǱY(�״I��<_�x��������:�5�]R�miR�IDņ7��p��a>ܚ��������[Yߧ=��=>]�>		,rx��8-�C�>^�����?%�B���d��}}�#"E�^���ޚ��O�V�~��x�{����m�f��!VR��`Ȕ�_u/����ؚ�z3΢m2!����t��������%?*�9ZLm�S8���d���j5�&��/Q^/�����9���j�?a����VS0�I6V�$�����DX���0K-���%|��Hy�o�W��� �-�R�5^��{"O��; ^�)��0b��=x��rQ�\}#䌻�rLGLv�T�w�$&gp��n������N]�@/��dn8�q��fp�t��qM�F~�]�+�w��q�$�&ۤ;xlg�Q�S3�����W㱭y��?�aD����N]O4���l��1�����.�O��q�B�\�I�8T�T�^��s 6n��k����M/�P5S�<��:��/����W��.%�ڬ"�I$2���$�z�%��7H�X�@I��#3|�2��g�8��Q4b���K<mZ��Ms�@ܞ�f#����]S����|⍗���̄�5�#}�L�1q|U�ѿ��-�Q����2$v��Z5�8m���dfGR�b���@E�Q~%s�� V�A�<o��)�����s���Wb�`�r��I�R�l�][j���O�Z%���ﰺ*�K��g[��{�Eӆɡ��l\Ɯ�YDãx�V���5a�� 7�/h�ͦD�\�������H��������&aV�ˠ��ۏ��S#��>�
�B�sx����!`p#�*1GG�m��F�YM�-��?�#oפp$�x۹K�����e�r^M`��>�&t(V���Tٞ�hFf��;�M���Y2�6�}��f<%�S�XB�+�vs,FuJ�+��
N#vcEr.l�cJ`�?髇(�J�˧6�r���?��͉�yЪ&��0�xy�<?=���	��2�?�8Q���]��^���.�O��2>k0���ra�C�wB�/f��
�.n�$�"��J`/�u�DNr��m��ݦ6��h�l���[(��h)�vA�`
�g��r8�?��Щ��@I�k�f=�E��]f�Z�Ց���7|��5�+t�PUCv�!�׌�u��ƾ��0�cn�����G�~
"U���̮ԙ�%6�e9��5�߾��c̯��Ô�����j�|��\�������t&�L�QKԧ�jf�|f�:yk/���.8�p�p����% #�/x�%�+�88#I1fB���Z�N5E%ސ�{��3�F5���K��ac#��ǉ��Ap�s�a����Z��"5�ȉ(���pn�{$A��`�C=͵G1�O�pR�.y� fl*9�D�3%��"������M��zʙ(������ͳ.2�c�y�_���F�lDm���"�+ɼ���X�[�6�&e�3�>���Mޕ�O�j��n�O������ m(�;qÇ����F�Q�}W��D�M��̂�l��ҒQ�0�}�id Q	/߂;�".;��Ex`�r����Ah|R��؃"���?��=\X3:M��+�W��0�/��%�Xܙ�w)�g%�Ǯ�{x��o޻r�~��a�A/�-�qY����<������r�MW�-�G�,���p�K��{�� ֬�+�7z���أc��U���g������2�f���ʚ*�lٓ|Jg4'1v��nhq��W{���g�(�kEWc啮���m���J��b-x)�\"��Q*�i&m.`^�����ľ��ew�L�}O51m<�Z�Ïi��:?R����|�� �m�V���D|��I ��p�@_0ѵ�}�襲-��I�EWs6tCА�@�
S�6,Q�G���?�W�[e�s�~F�pE}�2��G�X�፪J���ٹm�L�>�-��X�l	8	��9�KŝοQӫ/h���|��Xr6i�%���JB��|%!��Q�]φӬ-�	-^	�:���j^�2�Ko�{���Ge�'��#��u����D�'����>ڶ�Z6VV�T	IXb3�1z[|�ow����?��E�19����V�i�C��ᘐ��@������V(�����/���O��~�zb�E�x|ɟ�W�����u0��I���yFx�5>�W/Ф�'�TtA�KBi+2��	待��z��W`T����2(�W�,�[�@K�ޯ���R�F�1�`Y��2@��"#�>R!:ǔ�ڋ�L:��
�ƾ����Y	�% �hBl,�������)Q�ʩC�y���c�P�n���?m>�RsggV�L�tK�.!����������:mG�,C]𻁖-y���5E6���3��^9-.M�!>�aG��M�h[��R�17�l���"^|�..��ߞ`��z���n&*RL"L?|za~ )b˖J�y�]^ϓ�0U^��M���_��[z�Y��rgA��GR��ݬF��d�DS7�p��F��Ia#}�ǻhB�ǬҁG��VR���H�4O� hW� ����\�P�3�֖9�!gv�L�X7d;��Ft��҇���X��d�a
��؆�.Q�̡N�u�`�(>N�]_��僊F���W�E�M���`�ߖ���	��m��F	��S���e^��ZdzZ7l���x�0�tDW�J9��2T>�Q�'^f#����}f"�����x���DVB���/�֡��ŹC����8�\y��5�<�)��w��&4\Q�X�<We�5,]��Қ��3�&i!�H�L�E{����sbWxj �I"��:i��ƞ+L",�1��x�iC�Jb�ᕡwr��ؐg-�}�D�2��h�r�Y�qIM��b�9��*�-�Gsw�� ��y(�=-�4��A��s]C2�}L�P����9�ޒ5kU�+ة�w� ��E���1��E�12��e[�N|�,�WD���R��R�����	!r���h��࿘v��z��)���Q(:~��4-�JL��v�/�c��
P��G=�D�~K^�~�X��Ѿ@�¦��9_d�di��ʻ5�p�]�Iz�\���%��s����i�M/^]����_�Bd���ִ� q�Q������{W$"�g��3�譟��������lN�߲p$���/F���!&ϓ!]�N#wN'�UK�f����B�/�B��"�����7uY���2BR���0:i����"[����ڞˈ�|�%V������
}ԗB-�.]g�)b�.� ��=��F�L<v��/���jk������M�L�}H��T{��}���C���^��n�B�R�~�V���
�Pw�%D����/r߸y%~���Ș~q�e5oƑC�D"��88�]�G.��7�@c��{�dQ�>/ ��`��m$�G�J�����}�*W��C�7VξL{Zg�5 P�)�U�(Mh������u�1
d!���OZƳ��8�FVt#���#Y[����b�4���Y	�rj>�|�����d���Ȫ��Y;;�w����<)��f������Yc�h1[��eTW#s����ؙ}���� �����Q��I����������׸e�,xCD�]
�1�Ey��C����)J��ïT�+�Ϭ��=�i{�/�6�w��.�;Y{�bwB���N��.��p~��k)#�d�d�`�M��4����g���h�]�T�Z܊) ��U�̆�u�ť��OQ�B�3�Q0�Gg����8:8;x5M�?O�Y�7&K1갳��k�3Z�w��w_�Mٕ�Od��E�O���PBA�_�y�1:
�yE��m��M�zM]����Q���խ�����'z��H/�D� f��kA��h�~�"W�#�X���%44;�����x���{g�Id�^㊯�ɛ@��S�KD_f�:�|S��M�϶����;׭s�����MI!攐�Z_wFT�(yk�0�c��n$7�z���D��y0ib�t0$�O{:�F+���z;H�`��6�PPJQ�)�Z�S�,QD�¿xt��)9Cz~jdiŋv�HY� C5N�"g�WvU��Grx��R�%���c&H#`"Mh�/��+gp6t�t��u��}�	=m��b����,�Y`��=��!털1���F�0��!K_|S�=m���܏����@t���'V��K>�(�w ��ݾ)�Ra��~��Dcv"`� �IeR�E隍��D�1�ۛ�|\уg1R�8��#�ٙ@�Xe�.���sO8B�_��������dl��qo4�|Xx�T\y��7��8���`c�֌.�q�sL�~�hE��aV{
�VHJ�v��;���Jj���!ݡԞ��ĳ�P�If�>������b�i�C�&!i�nb��&਷�ANǵ�N'7z�z̸YL|~ajs�!��ff��P�\y�hb[����P�{D�M�,Ltcp�7�L��Zt��ڰ�U�����)��ұV�" ���� u�{�E\`��#�"�?Y��ߛ��?{X]��SVL����1F�@:��3\��ȝS�Y��|۱���Sm�+2�m�q���7��[�\Ey� Zw�����)��04 ��bB��m���z��}���8�$*���l��՚]D��ks�,`R	v��K�[�����^^.[�b-Q�w�]��g������]c�~yS}�j�sD�%Q�K���2�e�hm�Z�*Hvd%��BƆ#��$����CaCƲ0i��)� ���f)2�S� ���~*��#�R�����`� ���~<��g�� ��O0c@�Uh���p�˔��sэ,Z�uh��Oxj��S~��֧���w�`{zz�*I�k�� ��E$u���#V���tD,�9v�kİ����u�~ĎCRxK&�b�;fd��1�h�#hJۦ��c0-PՅx�S�E�3ܐJS��iBқo�"h�I>
l��_V� G��¹�J�;���`�@���2=l����T�Us���[W�שg�\��l:�z�F��҉�<�̾�+���7�uL�/$�G���r�U�uEH!��5Ef�
5�,�2V�4��y������-X�.E�J/&5�P;s�R�ݥcC{:�^�_�6���ّ�qq����G��5$L�|���Hd�w�gs_��ic��K'�LO��h֜�̸9S0�Lc�'�HU
6�'\h_�n7�ռ/c�å�gz1��&����}9�p�g��rzSu{*��u���o��fɨ���U���/ѐ&(�;����%=�[��"�. ٸH>��,�v��$�ԗ�Y>-S���g�m���ڴ�2!F�goyAQm�J[1��d��}M�V��ח��m$̧�A��m�]H�����p���������|�0<J*�o}er�,8��ш|'p��O!m�`�n/re\v�d?J�E��ޢ	�
��z<]gJ>Ò�� ���0g�
�GS�� �?�_������.N����(��`_s�^�#:>��b��eq�h��Z��L�Z��R�L�T���A��6X\�M��C�`�Ȥ�\��wvs�ڭ��Ȩ�9�_�����7W({~�9v�hƽ��F�� �����E���{����-��[N5Qnf����*������^}߈�
dK$\A�6!��,=� ��Vɠ���+�^��7����t��l�02�&"#~P){@z���DX�i���/L)G@�����WG���~t���ƕ����ܽ�c8����Ժ�$�#h�MJ셚�,O	i V����TX@��"��xŖ�X_	��t��PXۉ�c�og��t{W�T{'K
�D�{�Y!����o���ɡ��'��F�ߜ��B�D�ڹ��,�Ђ��I��v�F1@��^��dSg��)4���A�	� �rQ?�8�Tț�o�4
l#a���+����Z��y���]o���n�|m��}�6����NX`��Fb����#��kq���"c�!q�\.!p�29(��b.F=�v�^���V�����7JQ�ޟUE�He~í_�P���Ĥۓ��5�5�zZ��j��ܕ�GҗF7n��|K�.3��6.KL�BN��k+���c�I��۵E���;`�ѝ��`�i@���<���œ�VN­��^��M-�H*gz_���l�>���V�.���?,`��)Z�#��_Z�X[q�NO0
���	�NӞC!�<�d�|�7����p�m�����}�(smzg9VF�=�xL��v��ȹ�F#5�Y��X� �/!�����gwu��9o����������.
�&�!.p��G������/��]1�{dݠ��hn�)���o��*�J޴�>��wk�N՞wʓj$�ɯݾRwR�D�-���D����"40�	V�T�@�Qt>�3�{;�p
�V��֌�9��F G�1��/��i�_:�v1���C��p��+����}ax"�ž��Č��/�wl"?7Z�����<2"A�f"�?0��m�l��`���BO�_�Cah��{��}97X�����MuE��h����	�Q��� ��i&r�ΆK�FHs�+!����(� "7P�� �:m�Y�j��`Y/ҟ�
����%�W/ܭ(��A��ڀ�c-c�ٽ�9��C@�Ǽm BaC��.�A�P�;�Q����� 3����`$��[�!In�9zZ�ҙ"1�5�נ� �i���|�7�] �k�s�Ic��Ѽs��̤n�+]��
^d�g�^*���S�bl�
C�����S������4�%��£�ٓ�p��\���n%5WQ���!o�{�Tp�4�V�Ft�,�t!����b�K�u_�ͦ��Q}P	�am^�����w��ƣ����"z�0/�S-�V8�yG� I�?��Ҧ=��򉲹K�������_b9�Z#,A����uȴ�ɱ���|��T�Y��Al��!a������NR�������c�>�8�}Ye
�m5}��R,��ϝ�I�/�x���K�	/���J�(=���q�&��+��ذ�z�k!oRĶ�f�&k�/�]yť��ы��L���� Ic/���E��ۙ��������ť���cL��F+U��_.��'C~^v�;�NO߾ٕ�x��{��LҚ��Y��u�vJjLZm��A+���P:9�	���8
	�m��5����u)S^ߣ
{b\Y��DKӦ��_�x%8�+�0�U&�C,� ����I8ZЭY�X�(|��dN�>��ѳd*�VZ�~�R�Ӹ��<�����~��Ž({y�_L�C�N�B3J��
��0�eM*!r�s,�da�nɇo��}F<A��M������J[}��w�Q�.�W�vWyvãF�a��|�����"0̛�LN3.��$������V�e��g�9�'����� jk?AHc"�6��5������|N�3��`��J�މ��;�*�N��`x���	GA3#ӲK;�R�H���f�0�Lp���X0.�o*ũ���`��Q}kD�v�K�F����kjVGc����DX������3d$U&�uuZ����&K!1ݹ%�֡!���c|���嵐TGZ'O�ۚ���,�xZ�5π�t).��W�@qE��!�Aǧ_���\�:<��H6��|�.nL��c%9�1���4�e��[8	
D~J����2؀.�hoH��T�w��qֺO*����� :��Qzԝ��Ý�sZ'�pOS�(�DC��[��c�
j|!2:����G�J���'�ǉ2!MT6�;��	/F�/@Q��C_�E�gOQב<�]ڱ��C�mnQI��]���8'�i�B�R2]�D��fs��l��]�m�4��j�����G��#�A=$h@�9p��R
�[�͖I]#�����UM&UÚ�}U`�ԙh}6K++�ud �����+��u�Sŗf0�#S�3������x�m����/�ܯyYy�>ە�7���V��i*zMd�1ͤ�.��uiK�5"�Η�Z��;0[�ݬ�)��Ȅ�d-���V��F�=Xt=:D�f4����ng��R�sɤ&�q3���9�0�>��O�0�)p����c���yeDE�en$hs;�>?F����z�[v3�k�I�#z�7�E��l�3����_��@��?g�]����e����@�oъtD'b9{���&��wG�E)v2�+C���9��p'v�c����x]g$6��i�S n�v�c���W�� ��{��Pdp���qFE�4D*&��&� �mw��_p*���J!@MCN��s�l�U�q��sw%>MB�N�T�Dc��RMK���>7�L-)s� 9��M��<[�BO�d��B6��4���(V�IȆ>hL�D��w�$���ڤ~c${`>�ȸ�5K>��='��c��2�-�rFm�E���F0�S�����??lخב���I_\M�~��������N�KK��X3��	���T�''��$�+~_Sk<./�֔�+0�X���1h��p�Go�Sαϛ9�v|V��#�ʜ4�8ƹ��L��	��ڞ|��=˶��I������Z\�^\����`c��n7.u���մ4C�|��sV(��S5�D=>	1��W6l�!Ow?�����!_|f���,��ߠMckEv�"���/~Oi6 �	L������4��z�N��}\��)�L����E<�\<���+yk����{�am8��A�,h4ͷ��b`�N��b�����5
�.�V��b�B%���\��h���ZҜ �(�y��I0Y&�2���g�:����Y:D�6)��5n�N0]dW%/�4�C���A��	��Ѻ��T�ȁ�=��l�т5��9ޣ�J�~��^�mYk�+q�-��_����� cl������W+�:�ɮ[��ӡ�����h/�+�Yx�-D�s90;������;:\4��نđ٢ÿ�26{�c��?�b�-QW:���D��= ��.�DCX}+L��͑C��V�\�e푦�?0?���l��,����7�?�����8�A�8��$q{�?�τ�m� ���u�T'H]��G�>� H�3�_+����c%â�HG
q�0r7+c���#�ޒu��>O�S��#�g�qqZݑc�5�^W;n��d=K�1�%!؟��e6;�ɔy�[���"~��N4J�J�H����`� ?�&8���@~U��� �K�W���Z���J#��v�|��Y�xř��O�&����}��7S�E�]"��Yuc ^3?-F�����V�T�ၷ��|_聊1��䉲1G/�΄y�؏�b�\{]��w�]����K��kb�.P���;��%�;��̓�6k-�6W_]�r�t�_��^��I�i�����������&>ɯ�[*1Ҵ��2��g�����背�K��e�D��bM�ŕ_�:Pi��fwii�S���d��g1���}�cƐ�n,��un��?�̨��qk;���埫P�ĶC�Z}�XRP U�b��Y�ɿ�X"w��P� �̬0���z�ձ�nP��s����VQŐ�{2��_թ��"s�A�(�3��%eB�a�U|�*`�p�I�	m< 0���:�#;������X��_x���eDF����]���!Mc���e��G���up0��E��(�i�P�b��|o�}��Q������F
ciP�e�(1E