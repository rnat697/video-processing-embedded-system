��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh�%�v��⳵�JXH<b���m��3��'�C�ZoI�-�N��Σ=��˨v��Y��������5z� �c5O�4f�y��rtD��'��z0@U/�=���X��*^����	#���:�0�Zt6�/�3�&��Y8d6��f�v_9uU�
=O��9�@�6�[�����y߇X��˲<��o�����az�0�	Y7S���\3UГf�i�z���#J�� t��$ _wI����lV��xh�Ii��fIO�������a����4}ŭ
ڕډ����>-���P�k��d��O�뭙m�����JB{�L-,h�?ʵ�򜼁��7_�Uw҈3���BϏ����_`m�A-�hb+��,=o�_�utck�8�8�vZ:lw�P�{��$W�p%�[��A��\�T�
Q3�{`�E4\Q7Y4.���G^Y���N|��2Vgz����2Mu,��QV� �D���R�����˜�59C�h�d�����*A�-ƪ�8�K��s�\��!� ���2$��@òu������~ M�` ,�"'��L0"C���+@4�U���;���zj�w�|�v���
�VC#��������Ϗ_��Gi�$<ޑ�V�ɴH�ƴ��5~�m�Sj��KSd�[�4�#	7��-���Ӏ��H����2ٝ�q�-���I6ͮ\ɠW��iZ8��,�Cx�q�ucʀ��=��h�X�,��ѣcV�O>+�W9���ΛT��N�6i���
�(Y'�p��� ��y��uF<<ޝ��y������o��pX�O2VG�7
��T�p�J^�¸�Ք��Q���������cU�z4|�h����юdm�������sv�:���}��{�4���v�5�A�{��>�m��<��jO4Q�ӵ^d��$AQL��Idr���.F���:/$b�*��:
$�4Ϋř�)������؅�(��$N��6f���{I<�7��o��S]�k࿧���~��犺�^&3�Ḙf��@�����u��-�`9��������*{��}���@�w������t��n��N&���[�G�U8,4 Yb7#7rt s_�g��@��ݽ�)D��/ݾyN��8��[��j����)Q)n��#克*Z#|��l3J�쑔H�l��Oϐ�q+��B�y���c�GhS�Y���"��ԧxt�	b�Dذ��\Xw��I8���8�}Ƚ�%*gq�����N�Dm5�$����瘌���C˱^�ܹ%��c�	�/��:��
/�
{������0�4�A��~z��K�7t�b�6�	�du��f��(�<8=l-V"2�m������r�z\�j�_u&&w�<��ᄫ �a�0*k�H�FH�?���'$�~t�<�F�T'�f. ^q�0SW�<������@`+S�'�\2RZ@Z��s����!�C��=Sco�d&�	?�{�$=�!oƁ��h�7��Gk�TrV�dI�>�=�_h��O ʜ���z����|5�!��P��Љ�������4�������#ӦkQ*���/<ۇ.oot�f�^hx��:"���
���j�*�8(�����CȦ��sd�F����ם�j���$+"�5���Kb���$���A8���v�ҼN=�EM͝r�z��S��F�'�Pp*�!ruW��ͦ�
|��ނOXP�c�X{㦕�bJY8TT�����tyKUU4S�=��O�����<��%'_�\�����W]T�
(t���ZL�i�)B/ƭ++�Ĕ���&���-�9=�՞�M
���G�']���'��?��b=���@O��'UE���8P.-�P�7�	ftR��Bdd�m������E#�?xA�Ax_�s- �� 00�rO�;��R�M��I�ڗM,'�,�ʑ�Ub�)�c��*_�G8@�Q�ʸ
�
���ɋ�m����K�ga2�]f�NT;CTo[ z�/Rܦ����]�7z*�"��P $]��/pk�t5�?7a~���xUD��Z6�V����F���ˉN��(��U�>9�
������0��.���UHX�#���K4�w�A//���IN���xȉٵ\�4i��O�<�l�c_Dp�����(��q/��7m�S�"����w��ڽ����P�A�Flc,J��@U/�C�Q&�+��z�ףi޷᱕w�Eȝ�����h�24�"p�b}�M騫��4�+wE���}�(���a��dHL��))nz:�C
��9(�|��Z�k�}�p���_�5ίة80n��O��0T/�9 �	�6�B���<�
�i�z#�š�����x��Wċᙈ�_�� ��?
����4M&g�T0�	Ջ[L�ɝT�%�|�Q3����_!&�Ws���M�@�r��R(f=��i ��N_��'��$�_��/��ΟN5����g"�z��eժ���_����G ʄ���@���̸=!���p1��y�G�N��V>e�*��IxUb�oC����K�r}:xG^`|⋭���@B��
~eX���v+13e�x��:#R/��>�������oL��i�M�Y�x�E\��Ng�T����zx7N�A�	��]�c�&u�1p����b8AEJ�ɉB�p�|��iRN�kA�W��;H\?��t�^��I���.��?�b8� ����n>�ҵ�A̰;(w_�8w��cm�oy�\-�{X\~��q�,a��r�4�Ԭ��g���{�l0_0�pyZ��(n,(]��w	�:�Uj��o����o��y.��AC��;�4�[C]J��u���^�dE��ö��T�i:��T��:��5���7��6[�m�-g|��m+o��4�{E�|�f�K�"�+Ϻ�Jw��)7�]�j��,���M]�,+�A��Ǭl�5��<w��r�X~e�6����]�G�L����i�D��"v�Q�<��%�Q��gGݘ���apX<}��H���ߵ����Ɣ�#��2���BèBJ=���u2��B۹�u������2��a?�~���K��##��'�����,�s�z;���͒;�V�;�f�qu��ʜ4��jJ�vҪ�)��+eU?� ���3�f
�=��/����"eNI�BC*���l��/�:��}27`���%�䴱uܥHjq�~A����yO��x��Y�.�>�XWT[?�dI��٧��G�s@�S2�x}v�;�QT�V�ێ�J#���U����.��H��(�����+�D����`޲�(���n���
Ӈ��.�����0̌k��ă���i�;� 帆�)(O�9�w���٪���:I�k�Ip�����,`���B��"�0������|�1٢�o�2Ҹ���w�@�ke�3p��?�\JP0�`'��m<�J�Gr���j7&b�S�i](��m+�*v�u�e@�C
�i������;�>=8�ȁ�:�����֘g���pGx=0�G�`o
X4�Y����Rc�R���� =|�7���H�J������2�<�5���^4�gO�ƪeH��%@Рr�9~��eB���7=�����,�[��V3,�2s�L��,Fy��{Vͪ�{�M� �3�nה���'wS��mq�u7�|+��6��3x���Ўɦd_�~�l�D"���4�ӬI�ISހ7���Z~	�d�w�D�FY�j�H����p-
NJ����y�vl:�m�t��W��ۊH;�"���.+�`$��GvA���S��\�F������s�T��Ҫ�`v�3_'ܘ�5o�-0!�����ٿ�oi�V	Z-�[$ܥ@m����|"�D���R�;b�<�@��m�7�,s������R���2uՋ#J���p�iF )���Z'Q�ƪ9Y����`r�d60�c�B��錃�U��Q'�u~s���^��%7_�&f�O�iSJ��˲G��l�㱁?F�@6J�w(kD��2ϟK%��u��k�M����tq�[�NLf����=�Twa[d�ɜ/s���TS[�z��0��5}��Z�γPm!#z'�(A�2I��4�ܟ�c�_	Hh;y	/V���D��eH�a�JI�8+��ݷq/�賳���}�џ�m}���$7g����/G�!Ȼ&���<J��h����9�k��3�2����[��?�]�=7}[�c��gWҿ������*�Q��0��'���
���|TDO�r�w�E�摔,���7��Ob
�\��⭾�����IoR +lIfNuJ�Ƹ>ק+���y閛WەR��U�}��)�*l��x�>Fd��E�,���Շ7��9���õ{��v}�9�.��-� f~����F%M�dr3��ʲ����"�/�@%�^?�b���=��
�x�_��`�OyZs����jpW�O6r���=�Gc���EL������8(\��ª��@�f�|�U�&���}�Z�V �@ QXm��� ���m[+NCiVϻ�߆c�	���ba�3iJȰא1T���>�m(��;�������v���0��֯(>F�"�X�
y������s�)H<�kvm��������E�Q�F��#OY^������/flo�������+Z�"U5�!b�+�e�9T�O����K�]`�?z3w.Nj�+<�������O�xZ�f�M�����L�����@-��G���v���ۣ�]�Ͳ���TLJ�C��~�O���z��1�7D��������	�^!����������%A�0���sfG���?������L�S%FQh2����B���J�e��̫��l�Т���w<���<��Ms��VbRK�1�1Z��2[o��$���d�C� a�(�zPfNB	�;@B��q���o�5��O��o/��>;-��r����z���6��~}��8�O��h�}��>�;mo�N�5�&b4#D$�M���Y���t�ę�DB� |8Yy81��H�a�{����#lW���Ɂ\�[�	%;j��T����*L�O�Wj��l��A�Ԫ�U�_�ܗb�M����:B�>������2�G�^Q#��T"�d�����7��3����>��~
��Yd;��rE�c���A?�8��ד��ʲtκ��i���N��z�9��f�1T��ցS�ke�z�~�kުM�F�ȽY���n�j�
@�E�iNHu�r��V���5�-�H�)|M��ZSIe���&�������� �'��J�v�Q�* ���I/��X�d��v�p���6�s�/D�9��D{��p�(��L*�
̢2�G��8��(2�m������K?�6Y�kd8�w�X�����[ax?���R�yA�Vc���b�/�~ۈ{�ݟ�s���]��������f�Ԣ�4�]����U&��S\����u�{�M!M�fs��O��� ��XYF7y��E�e��5��׬�@G�5>�0C.��57P�N-y��X����sN�S*��`�Lű�X�<2����1E�M��/�`c�<X�R�7Q�h�n�_��e�9���8>�f���5,�;���i��F�{�n`'H��^VC�K�"&Aׁ.	�*�<g��Pj� ���ko��hs�O�%����&Fcb�	
�:����X��n���S��B*4�x�B�v6�DM���e
�m���m��3�u��χH�(VHɘ���{$��a?+qΊ�u�NB�������>�|��=�z��>��E%�����Wo`5	`1N�RB�E�z�x���A�)*e�LH���z`x��m��R��9u@�Շ��]�>Zz�7Fl�+��I�4@O��D����V��3���z�0�t�U�S���r䠎���h7~�f5G:�?�1!/�9��er4.�C)�*9y��L�d.����?��{��ݣ�6[�)K$��[��"��C:c�m�/���N7�����3�v/�N�f{n�f�x6��i�7jAl��KvZ�U��.��gi$	r��v�����z�R��q3�����6��{4��{5����n���� 'p���'�ͮ\�l���*S�B?�|z�g��:S9����V0Z���l+��r�ͻ�b}�Z�d�00��@��h����k��Q�{Lz9��Ӂ�[��]���{��@��+Oݰ��a��v��W�z�O�Y�[{QB
[[<���b25	�\jiB�N��_Flh(��Ψ�����I|s�OEF�H K�^�*�!lSp��fi�s-�#rS�-�Blk?����<��B��!yD�Vf;�Z�G�SM	~`)~'�+�����i2	O�"����Ǔ/�3a"�[�ˊJt#���͡��A'�����DJ}�HILWxL�#W췑�Z`x�k鯈��[Eᓿ� �Z� �GG���2v�!�m��v�-�C��9<�w���qx��>�
 �-A��H�{�x���J�Nl ~m���y#C	a��0��A_Z��q�)Hrt�����8e��rWEqg=m��	�B��țB�\�T������[��T��@-`��y�Fb?I�i��>�#�QH��.�7�)��H۾"0��j\<.X3���U�Aʣ�6���.%�?؃�a!����#�1�_�g��4T"K�N�8\��Ej�p2�W-���a�V���F�ŗ��^cL6����<�`)�����6�)��"�*��Y2V,�)AAU�~���Xメ��s�%^(g�1vQ�-�W�8��3j�7h�R5s��^'ֹL����e���`{�M4�u%������ |@&.p�Ɗ̙�c�"u�,l��ell��>�P�#�Z1���g��I��Lr,�E��uc��G�p�v<O2�u��"�՛|1"�v;���k�P�I��q0��	ݣa/�����z����@
�u�c��][�Xʍ��3CS�f醙P�q�_EB��2�/�5�o�fd/ji8��PIr%{��Y4(��hn���PT)�mw�˝0�*�o::T/�Y7�{_�=�,QS��&P� ���v��E�5/�ߴ^�UⱻQϣp)��s��Y�[��&��7ͅ�5=���\��%���ah- B�s"x9Ӛg�v�h8e�ʹ���q�b{-u閱5VQ��cV�9^|s,�Oj�E�F�E�5����|�ݖN�>LW.�n�Z��WC����"g��HP��!�%� WQ��񡲙�iv
E���	����F��Gs����4W��	�7H[�u�w1����v_=��ç%7w����c.�L��m�۫.fSi}|{�h�3M]�%����?��n��T��&6�Xp��Íc�W��5�,GqzC���C!���F� ,�4�z�~Tٺe���r&��Ɗ@�j�y�՛|�j|���\"��WQ�`I��2����{U�]y�l	�K���w[گ��l���Z�����ȉ<f�6w���Q���RJ�S�q�
㪦}m�(x�J��S��G�ُ�s�BAj��E�����3�#U�+�B�k�r��擄K����b������fR�w���S�	5���&�[��Lh�Ql}�%�RG�̵犸e�4�˪�aO�S�+��Bozn�2��e�ú��X�;d�����<>ucq��nuE�a�Y�)����mr�h����l߽��Z�g�cx[�^���Y�n�d��#�VGdg_|�K9b =�B�
��j݄g燞�,��<����s{���Z�H�|��{��ʝ��� A��qz���)��G��CM�Yb>�a�o�s�����L�j��S�ă��j�lK��B�VUe X���"ʬ�h9���셦���#p)[-�bP?�`��B��hdA�E%⥮W�F�=�q-��-��
JtwB���{���o� ����yS��t�k���K�)�%��c�E�}TjS1��̅�y�b����:��O��AaM�qjC��=ͼt�<�����"��k��+0�r(*ʉ���U�'""x�ݴW�I:I�05�6���d���[q�@P)j���/��)[ζ�&n�Y�<l�89LS7�T� U�frЄ9�W1X�5
��IC Kɯ���<G�Bl�z&�����N|�&p����R����Le�PO��:����gceȢi���"\;_hC9Fn�t	��/c��_�N���up�2B��	��hj@��LB_�{D��Βo�|u�wԹD��!��~%��(A��(L�-�x�,U�
_��{�F4���\��Щ��4���SV���M"���߄Q�$<�?�|�\�|�{�nK���l���؃�+�i��Ȳ�+˚E@�5��w�l���n�cN�'k�Iy;��/?�Nu��d��\��v�R�H��/�+|�b��\��UcD�jO͎q�[�3���o�n�T�����
 �XC�(��L&rԷm��k��o�k�#��W�,����8Y��?�D{�_`��(7zT�d[�w��Q�D]�nhA���&e� 8��H�Pn��߾ �����,�3
$\=9��y[Q!x��TK�!��dW�۞��k�R�v�ˀ6��筳�қ_h�Y^�\=�b_A�����ڥ�U���l���</��|M�=�x�{�1�S��
x�F�:�A�>�։�a�0��
Sl��O���b���Ǩ(ڼ9r��A�@x����W�L�0
GV����g��E=��'�Da���"[�ݿ/�dT�����
�Z
' 
*K� 2�Н��*2�_�̻�H/�]�����4��L53^!s�!̋Z�É�^Һ���ɀ{�߄�2��,*A���aUz�v�ٿ��@�[��� _Lo�cͶ��J;�Aw���i��Գ$�,E�ع
L���^��Um9���k 3��fO{�8���s���*�0m2�e�6eO3A%�� ,�yd���[�L�gGS
)�"�*���<�$O��!D������yŗ��u׼�dS=~a�h�j�a��J��/��u��+�<�Xp?7�Hv'��{)����e�$�z����튂+`L[���1�7��)fׯPoN9���l�^^���@	4�F��/b�� .�c��&s���BI���.�*)#�鈢fd+���"i[{e�ܤP<IM�b�(W�iPD���Z�[i�` ��̉�nK�ɧdo<���&�"(#,�o�����b?i��n9Z�<�mAxk�<���7�h��*K�$$8 �hY�/m��~�M�#�M��#��i���/e� �4P�)�.�<L3
�TL,����u�X\�U
�z�+�p1�� �_�Xe���d�Չ|�0��{V�[qixI� �M^�����=D�e�R�'I�
��WЮ���_\�\6�b�����Q�Tj��d�邒�^E����\��K��G��c!�&��x��G�dj�x �$�d�����p����������\ێ1�@�����St�97���8��!�5q�ds�pC^�+��9Hӣ�26��+�^�d3G��o`�aُ|����>�R���RJ�$�E����}�N0�YFͩ��h���A�n��PY)�I2��rX@B��/-�Dx����㡋U'd�1Iݕ�&�c9cU��m��egCY���6}�̀�Hv�4ŧ���sHG'X�t�=����J���{�2�EGN�=�[��KX[kF/*ك���'�D�g��OIZ����f�e�fD��m�G��>y.zT��v� �b=�Ԉy�/�=8�`��L�|���p��(i��z��hB��V���F�C�Hd�^w�	�OA\O��H�N��,e�����i����N�0�fE�*�:�SexN����8z�S7���UhDb4oNG���_�C>��mPG�,y~�V�g�l���75�(ʏ�x՟%k ���J/VE�JE�b��.��.���h]�R�
lވ��DN_Q�Î��k�S.���#\ٵ��3��M3��Mi(w>v(1�0����9p�*�$S���t5;@OK�m�E�����BH�t��\�xC���ٝ��ͤ����%j??�������$�[�;]!��r_>��V8g&�H�������}������L蛕��I�������ܡȘ��Ie�22�0���1�<%�J���Ud�x���4�/�c�Ń������5z2ʭzGSe'��M����gX&�Jk�� ��!y��
9�$�#�g�{"��ܲ�4��ƚYyu��n����9������Na��;����ݞv�_1�c�ς�˘�{�P�7���dZ�WΜ���6�hUc�&�����P�_ LD���N���/v%��/;��k�Lcf-a;�/8Y��s�����SpH�u��I*�Y�H�X:5�D�'�~~O!f���#��� �jD��&�&��s\�4��	��L�.�;�*#���ވ	���PtI����mlwF�f֩jݦB)U�=~��"KqX7�|��7�1��DU���D��˸��D�PY��h!HΧ���I��(?�W�x���n|o�!{�;9�)��H��� �b��¹<�XK�/�%1S��%86{#AI��(w�gLS5:�ֵ(%��s�����1�I�c��-YD��B˂t�-� �u8m!}�����ev����%ڂ���~%`��[�P�hq�n���ǰ7R�+�Xw��BJ/X�0S�-�����v��q�۪�C&M�Zdᆷ٣%�|KXz���Qؿ�:C�ԛu�A� �J��<���G�}D�/^_��U��M໥��}p��zz|1���(�N�gc�i�ܷx��������cwư�n��2���}�ʾz�0�*�w1�m��� ��E��4@�>�l��k�/}^�I`���wh�ד� @��*�qe���c�	A:�ݮ��4iH�b�MU�Pb
d-ؚ�oh�[R���(�W����v\���y
����;Z����ml�}<&���$Լ��@'�s� ��@�2��l�[θ��ƕ�z��{{v~wQ�5x�l&�xR�]�_���C�2F�)��h#�	�*D�1���W[�Jhlr��t�=G����X�+�zs^J6wg^����x�G	b��U#P��fN�j�d)�Z��7X�� �V���k��R@7U�%t��=H�=��;,�A&��&��׼c��3��ҡ�U��:Ȱ�~q����Bc� �B)�I��.p����	�n�jj� ����#]G�H0�g����i1�eȐ|[0E�>y��`]�r�}h��E!ٶ���Ul�+u����� [�v�	mH�F�J�<�Y� b5�[Ă��`�( �GN}��}u8���>��b;�jma�v��hp��n��t9�Q�u$�'���'�
qo��ث�'���	4�@�Ք[�f�!AQ�Z]��%����A��l׈��U�Y������Օi��z?�ߝ�:����B�p*ð��Zr�t�A�qR�-ݿ(6����_b%�Z���֯6��4��@z��m�~?�G��������j9Rg������J���<����ʤM|5ɄGƿ˛,K��bx����'���m��p͒o����s=�-��ʡd���(s��@},���\�h@�z]��h�Ob���n���o��ht2!��/P ��ѝ��9T�%N k�7�?�����r�K�\��BۡJ1p�ߖi>G�n`kF�7�v�E��m���k����T��a˦F�	u�C1�8x/�|a�+����k�U]JO_߅ֿ�ޜ�����ׯ����z�|E���Op��	)wW��)j��N�I>_��Y_2���a�U,Ɗ�L23-�0�C t�qF���Ի� x���⨘6��8x�O���9��c�3�ڮ����ZE��X�L{�N���g;?��k��e��,����E6�B��[�9��Y�W0}�h�X�	ɶܟ]�o;�����Ob�[��>nM��d�%��u:e���>��d�%t�y"y��
�����I���g��y�[8o����{'J�}7�h6�8����������J�S���w�ؠ�����}�f�"R�E�8ڂt�#i����t�j{�@�=�J�u�@1����s��QZC�dΊ�lo�=g<C�o�1j�œ<?�%��I��_6Y���x1�!Y}^�xw�Tӝ?�\�-vxӏ=�h�p?�� %Yi=Bj)���J[��7�������<�r�؂�����
�yUJ�NTc��y�f��c�q�g�:Nr���#�eȐ"3�q�q���5�7��_��3P%K	+��g�$�{@=�wh[���AbR��A#L��*0�F�����m�~�x/����q�k������	Xs�j��A{�I�/��"���h���U�8�&W]$�P�B�6���^�dW��1�p���X�.3Y���N(̝�iM�g�b��_4��z�J���a��3J���_���qgʎBF��fB�!�Eeu9CHo�"~�52�	� S����M��Y��[�4Xg����%�ܹ�G�"�Ma7�C�$�D�l��ĺ.�?y���_d��m��n�������i�0��o/M���7�OSڝ#���WP�͙�U#o��G�hM�Fڸ�/��CҞ�n�<��BK�%����5b}�Q}��spCRRc� Ε�{M0����fny��`gTq_ɒ!i��0,a~F �����U	(�|+:�ѿ���VM�qZ��\5C�sw�վt��uN���B�B2�w�Z����L�%��	uX�c�gQ���t��>�aw��#Մ������̵p\����"��nm��|ĵ!赚S��{�=b� �y���;�L G�<`�sdE����^�y�y�c������N��LD�I�������V���z�� �3�6��0dDZ�CZ�L�7L$�\y$[~��779~�f�DiM'��A7����d_�Y/��Y+&P4�s�˜A�NL�(6m�����T�Ţ��z�`��<��">e�㤚q(~.dc������l��}d��#��'�S��䜢�҄k�%i�H��n��Q���̟��v�E��5�(Y���S:���@HX�Z��%��L��S�js�yo�y]0Z{����A	n?xC�Gt�V��CS���İ������pd��[����%�]����!8}	�u|�{�mu��Ȭ�- S����&�a�I�G@ȼ
��4����H\�~�g�IS	��E��Ba/̫�j�٠�����%�kh�؉K�
h���	3
�hHd{y�v�_��zj2�"��kHc���ᛃ{����E ��-�1�0O>i�����W�#�4]v���v�-�~��,�ݿ�O�xƚ ����u��aLE�����I�#�r^G�����h�*v
KD\j�j.~�]���R�<[yo#���^�w�қ�z��W�\��\>F�^S� ^B%'����.'ɺ4�*b���EC�o�}Sv:��Պ��{�M�}��	�K���E	�|�i�ħE��ȓ?p����An��`��h��6ÒW)��.-�e��Բ�1qk���:��GI��pE�s�/�� PoS{�GyU_	c�د������7b�͹F
p�����X��"u���>5_r+�4��c���C���A,eJ���V� 7�8.n�@�ӛ0]���
O�x��G^6Ӳ��� �� O�R(�C�z�/f��)b��RG����hp8�!�p�8l|(�ΐq����A�-Z�#��O2H0X��o=h��dv��� G��wۨ�1��_�;��Јt+!��⽷�����^t#��\�Z��Ѻ�51qV�����Vs�,>ԧ�kw�&K#c�D:S_�e։�)��9h��fՊѣv؝6M�cq
?2���@��#3[DʐZH{	k�b�d���c�;�"���M�	d8��I_��H�~�'7���H����9����P�`�C�����譒s�:i��}�����c�xb�y�SZ(h�?�G�$�^�3\�Y\�W� ��1q��\�� E��	!�H~L�d�-���<�Ĺ-�|�e� &�����w3�t��gz�"��q�TOE�MSsa�e|��︡Nym�<�Ϥ����"ٿ��8�J�v=������P ����9���i���*ޢ@E����XtulF�!1�f�Tq����^@�9�[�ZȣM�4�����@K���D�m�0z10��1�v:y%�Y������ڜ�5��Jդ��/��R�S�[`�dmX:}Y���a�hd�#+��va��3[`�=:�'�u/�1�7�����O��u}ಔ���(��O��a���]k�v�{�ց�/���&��v������2���M,x��V.���R��I�Du�)�<���oA3&����K���Kgƪ����N���y�N�n�zDy�T��lSq�P6#j���\{�*V����/�Y�M&3?>�/��k_=5��.�wC��;�ުϐE$� W�O�d0��E�X?��J��������) ��T���5�+a�}��c^j�~H���@����dNs{�^s��D�b�Х�&o����pbT���\�{����b��cwrff"�7��4��\�M�^֨� ��e��H���@�h�~G��{���﷢�A@rț$��4�A�_����~i|뻀HP$3�Q^[kSX�N6	�d�>w�Z�����gJ��dl�ԅ
 �=��n�������\uwð�ov=)��r|K�(�R���l�E����v�4�=��`)�Y�A�X@�?{�5^t�c�����Z��^�m���콩�*ApP���#�c�$!=,�6/s3QƱ�Z���5K�r*�j��}�CKcA'��(c1�(da86+g"�e6ԣ%ż��zۻ����6}�]�,���Z�],A���b�_��\9%�ʼu9v���JT�W����\�C���4��4��Ɛ]c��u0G��2H���OW���ꏸ�z����A��v�m�cơ�1������'�����r-�4z���ǎԴ�p�M�I��2�"xtĲK3\�<bŬß:ձ�zH�	W�d��J����ci�!A�j�+Sؾ�L�5X(�V �L�?;B��d�I\*���ױ:z��߀�Ng�9C��F���1T�<9�!�R�Ju@v��x�d4��N���؁��_���O�+!2/fN'��1�KY7%�����KVr6먦֋�$PT$ ��w��1L�G2o@JE��Y�i�[��TC��L�	<N[^���;�tU�;���z
�"��s�-"�b��4+�Wm����ћ�rT�5g�����r�<c�#�������d��O'�;}=x�1�F�Ē����^���_� �)��T�..�=��$�<FV�����;����#�7^�o�;ɪ�6(Cβ1[vz�P�A���G�2g��[��� L=zX����)N7Ǽ0rt�֤m�