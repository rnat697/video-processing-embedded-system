��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�F����c8�@S�B���Y�iO��!W#��,��r�.��b��%����2m��ܛ'�*��1��Xq�U�g �?�8`����i���q�y����k�8r	�3�\Uz#��\�R~��+?��m�G�)��9&Z��]tY�X�1I�I�]We��8�~Gu��O�;��Q|ya����v���t���uZ��(fcf",ƃ�s�3-� �DE�<l�s��vN�¦�*���pJ����ݫ��d\E��d46�B_�Ub��΅%��>���,�JPnAt���{���n�9?,��*�8��izF�㰠|����O!Y�,U)i�{`:%�do^�*1�[�j�0@S���%�X��)
�r����/i���|+�]B�~+]����i�R��L|�����#{��ń���@c���'б��_��X$�a�t<.�����ئ�^��W����6�>z]R�E@�N�>?�P��3�r.&Hj�&�aI�3P�j^����1`���؞M�L���Z���ڎ���|a�����䎔�A���Ɂ��`v9��S�xJD�P"�v;�p� 
�%)\��y%mIβ�}�ٿ.dz;
��x�������M�7��*�����ԵE��pS�ǹf��>`/R��_[�b� ��6�}Ɵ��]��s��MӃ_$��kѿ����7L@�[������Z���: ��ɑ��n�v�_VY!���a{h���ր&~�O���̿�x����F~�ä�n��.<q��e�˫;�c�����#����zV��ni)�\R�Rz{��]�B�Z�i)ӿ��:�s�ߩE$ӕ��-���m�;|4$d��P�.��v�#�5�q��WсAl5�����ç�x8/(�^�K��؃Q��h�]0�����T�����%�~���g�J��� ���Y����`uiA��7���h� ����\�F�����Q��(&���G��Л��O.�4�? ��>G��n_ߚ?���FZGjYź�H�gޘf�3�'��x���7�h���#CA�U�!<&� z@�,��Yhg�PK<�C�P%p�&�i�\�׿�3��pe�MkZ�h���CI4�����NH
4��T�Ԏ�����eQ2�)�O��'5V��o?�Ff�t~M���
�=�y]J�O%:�+ޙ��8?5j����o�i�x�9d�T���s��S|���� 3 ���G���pD���?�u�# �p)��~y�+�s�jkH��/7�"�EO�*T�"2as��Pm�̖�h��v+�4y�n��|�s,a�,����+x����P�p�n� 6��V�^��GHk��z�L�^����H�&�ݕ㒻uZ����Į�{鳺R��#�Z*܎5��U)vbI�7���t�Q��恅�^F��-N�Y*S�ߦE"~��y�T�JLK�g��g������]e���YU�*v�5:�d�J��wX��E�Y�W<��!!H�?��¢���&ߟ��p�D��,-'V~A�ÜK�:�V
rA�dܫ��Br�-jR�N�@|���X��^�;B�-a�JM��vr|K��+����c"�ڑ�kۙO)�e����d�4�����k�t3o�m�`LBr�/������т��#��`os���e���*㑍n# Q��<�ԆJ�X���6�6(���~ l���$�~���)!� qNp�E�n/��Zָ)j3��a����
&3��13а�1P��ى�Ɯ��ǖN5+ ��2a��L��
���լ�&�I�@��b��zi��W�֥p ��b�k����Oh��&���#�\?�cc��N��Xd�^�>-X9�7N��j��կC$��
��}P��^�|�^�?~.�aE��*r�q���3sݩ�E�Zrgd��6&����j�p��U�RY�X�^Ⱦ�X?J��O�<��6b���� �د��9�\b�fq�Xw�WJ�����WW��N��*¥����b
�@��������U#Fo
2�:�3�����<57���}J܊_�^FpM߫!�L���H��5���h�f9�:x�pQ���8�%�E�\BH3/,S0w�g�Q��� s�Q5��f"�M�C��]����g�b��H����(��ibUN���q���R_`yQjK�f�y�x�	�^p�F�}֙�������d�J��t�[�Ԓ"!Z@|]�$h���?<��� ې��V,��v�\����ճΜsV�f~&�xk��BT�8{@�m�kY}��w鑊�D����#�\��Y���ĳE���ܬ���ơ��-�A���a�i�|$��M��L�[�Ə��8�,u���'��6o�x)$A���۾����|H�c��U��M@�0`�5�'R4X�]��-սM��c���"��KaZ'�T��C�q\t���*L����D3(���QYvDc+�*��~P+*��i��^����䕊Krz�� Ū|_���Oϣ���m��T�A��N�w�n�sC��Yh�����ό�9"nyzd)U�G)/�Z���)�ףܕ����[@}�߳��:;$�o�1�P�Q}[�)W�)4՛H���*���v��d	��иh��>D'cA��My�k�B2]��RX�Fё�P`}�]>JdWsA!�b��?f=Ѓr�����%�>O�n)�|pJ��2J�����$�D�� ]!����m�c\��']U�7�30-a�j�e�0t�L��%�)l��.��Ɛ�N�a�	M�*�� �J���?�#O�8�wi ��D��@|ӻ'/q���WusQ���b$��2�m����vҕ۳�ƝGl��⸫]-�C���5�L�����Q5��swN@Ά�E����\�(9��ڇM�^�\��Hن��g�#��=O��
��f��u\9lPJA�~�1�Ъ�.fxwE���p���$t�p���SH9�l :�5���yJ�͛H>�\||/���ީ���s+�]9s( 8kU�����z��x�q,	8��(@�i(�@����a�qrK�V/쬏	�oJ7�����}U�'H�j�<� O�?�eqj�k�^��`[��F7L���d�i�T�gn2֡�6���t�Z_�!c!����9��靁t9�tC��}]����ڙM�*=f`d���fR�`,6�%�2��a%_h�y�%Zw��@? ��6J����3>�@84��h�E4���Z`U��dH!B�T�t�df���ĔE��9�0^�}Jw�r�c���ٌ2�<`���N�D�J��I�Iڰs���$����}0�\�n��X��о~j��8B���[�p/=�<�9\��C�1��Yp��z��gf�чu	��TO��}P0?�ݲ#���Qi��D���t�!-�<�}f�K�(��'j����%�l0���E�싖�Vէ�����x�,���[�߄c��v�_Eކ��i�vj
�P-����W����f��+�
}e5V�-�C���t˟�)���#�j�ٮb r������8��v[������:YfYƊ��ruڙ*�������&\G���u"稚}e������O�8�)�����
m諍��s��������n��}JEF��S�{�;}�b��seH�@-9�R�C�P��B�AXgH:����|;�t�D	v%s�.g��Lg�?0�nμ!���;�E^s:7�l�A`s��ԴwQ���.����33=xK��h�$_	%���~v�[� 5#0")���߽�1Nz�?A������x���W[��k��Ѩ9���T�O�	����:p�@��vy��(�qZ��{�������gU�[�G4Ȟ
0/Ѻd�i�-��jЦ��M���O��X�;D ?,�����jȱ����`�X�3wVITFɕw�&p�R*0���~���ۿ��φ\?�zT���#���9YV4�8�d\�9�$i�f�;��Z��tDw�X��i�1(�j�0�<O�f[��j��d꺎�x"p-Aw�Dp�,:��R�$0�����&�-G>N��\����9���m�\6��Ρ�O;KX�W�#z��ū߄_�+�д}k����s�,����&|�l����5nPWS=�ܔl-Gi&ԫ���TO�u(_&�R�`V�D�� #pv���a-$��A�O���B?\7b&�9��h��nE��F���|�@W��G����5��в��VH"��5�L���:�N��[M��uai�ZSJ5W#��Ć�*T>�5�l����~xU��/a�$���7 �v���A��^N��uBH�ߴ�F-&&��K��8���/�+Mh���wT�A�vq,��YO� s�H��V����w���8\D���ʣ6�Ǥ2}~/�un�K�k~��P���W���~��B˼�P���$�4���%#���~,m��G����zT=�Hc�/f%̤}cA\�O�H\9��5��r`z���61�����������?���V��ԣa���j] eo���{��]5��U&�)�p%��^N�1�3��XH.���{�T���4���0���C��>���j������o���+!�и�T�3~�U��>Ϟ�\�PU1W>���Nj}x�d�/�O4֘����B����By6�=hw�H|��=2�zt�|�k��*�9����|�U���Ώ1���Y�GC���B0SJ������{n>�$�$*��6��Hf-�0E0?���W���Y��LpWT�JM�ccB��v��Bl4����]*h(6��G:SY"%T���Z�ф��3씣u�b]�aJ����;���W��I���Z��N��N��3�B��n�ß�=�`�x�P���R�@��kw<V�?���D�S��(hD
�D��KW�����"bO�-��`�ռ?�K��7p���21S/7c��ě@#�:�bw��N�ᰑ�������w�1X���-�/r���RKUI�^ �7��Y�y^|Y����H#��T?"ᠶ�Q�8�ڎ�/���(5_נ���G�ϰ�c�i�^M��@a���|����.}�ˠy"�⮁9�aYR�<�����KnL��L���F'�����Z0F���2:��:@#���D���g�K��7WK��<�{.�4��n�h����<3�M�C�E?�;�}�~0B�F�'@�BϽꋔ�#;�(�ʔ�N���12 4��7�::1NયjU(�����#��]լj!�|.Fj/�g��n!���N��">Vxv� ��v.хy��ݬ̫]���[�?뒙����IsN�$���r�v��o�S��wnx�����0�D	:oŠD�������v��c.i���>&��8�J�DQv�i#��(���ߣtl�"�?�rYql�4�#���L�L�"p��4�>�7���ܖ�6{��U�ǦfR'5��^tЧ�[̙��AbB��B��S�Y�d�b9L궩~����:QLoΆ��l�=w4p�fJ%��Zد'�v���䤏��U-��%��A:d&�JK��v�,����=!�.A�E��<��@j.(���a!Nu�b1�=����]��iıN�2�|����W{����Ǹ��{�0���Z��.thg�"pt��Λ�=)sD�w����( ����L^28G���\qjRJ�SǬ�8i�H�R�Y�X��>�z�x�!�����Z�UaB�@��t���h�*C��c�2��r`1^s4����=����(al�W�"�O���?'|�:��;�����ق��	<sj�}S��+�%Ö�1�1Оo�x��x�ή��_�lLAO��f��}�h�L��٢}!��VE�5F���6vc�Wug�O��}-���E�3|Í�M�a��1B�f.`��Z���x~��Shp�G��D-��h8K�{������Ը���x��v�ip��b@f�e���L��Yu���0Aڹ8+��r�[�65��?�缋�%%�P�6q!�~�Rŉ��
��^eE �(�y꫎����H� ���Έ9�j��%�� ��r:�}�h�~�"�f��7T���ߑ������~�q�g�[�9b�+b�Vj�yB0�v$d�؀z^)+����&�Fa�*9ra�c�]^�d�;��Iӕr=ф�\��m!I<�>�&��}�����w����yD��ٿÀ��6=u1�e��b|Q���B��ɛ")�8p��ꄟ�B�OD�G8=#ݮ�[��:պQ|B5�_(n��A��	�uH��pUA����]ӈp/D���D�]�ӥ��ԍʩW4 �)����F�"|�;[�t�/���S�ww���`��\�������������B�MYC"��=���F~��(��+e$���u���|ZV�X)��G�z�.���]������ۍ���{:�x0��x�l��_��)�L>� ��c�&T�c\�T��e#���`$�C�O��ސ��6'�P���M7�Y�֬��@|���*F(;U���AS�z����
�љ�{gK;���!"d�Ek"�X/����> ���˙��Q9*(��:�:�QH6a٘'iק��B��!�vF�ì���$��P�//�y�&V��j$����e�����,E�B��[ o껇)��vs'*����Ռ�aʅ	�V�g9�2:E<@X)Eʰw�!�g0|�����p�~]��R���ud$�$���ٲ�q	��\uX>�u�B�) z���6M͛z������/%I6�w��P���,��.���9 DX�4���7�Iu��?���#��]C�W��,u��el�-7���z{%��#߂g�Z���}�l��̦M��2����dlIh���cn˺Tge�H�p��=gE$�����wE'�������D:&)f��6�4m��W��FR�G:��S�K8��=�\uK돣.�R{ƚ'mw`	K�ħ��#~v������|0�-�^"��D�]��_V�^��$�%�*���͖K�k��ӣ8S� dH�λ)��%)>%#�x=�r�bl�S~Ы5����7�J�V�"�-�)��P#����&��,�j�we&[\����BA��R%lƔ"R�(�ޯES��˗)�>����]�-�X����u�����J8�{�O�<�2�o:V��5�!Z�=]t���ē�h�0��}�s^�B������Ÿb�C����DNf��mO�a��&}���F�|ՅY
c�oL�����|�L����T+l����u�s?�,0"f��^�r1T�fzi�L���]%ݟ�+&l�i+M���Ol���È�i8~Tsw��]��}ڏ�,�dD�^����	�A������"�MZ=C�p2|[mK��� ���Ӫ��G�C:�d&9��G$%f]���V�h�y[���Q��OH�m����񵸃t6�YnZa!�(�����K�uFt���`EMދ��m�[� �N#�v�:q�ϝ3�����P�e;(�,}
��4�2K>�9�z$lZB��i[�o	�fI��\5ҳ]ҽ�S��7��S�<�� �ю�D�f�d����Ъ��Zvwq�C9�lcM�y����;�)�Ŝ�B$�n k��)�W�J��&���˓$Tfl��5nI���^Q#�x$�|�e�ӡX�'_5�I�78!p��'�φ8)PC��O�&J���r���+�W'/.Z>�b�	o�T{�N����?�v�ǰÔuxalA�b���Y�Y���~k��rYe?�z;�8�ʇY-�c��D�4+�}.� �N�a	0 ���1�r��;��w��� X�E���#>X�a����r	1�[��y�C~���N/��L�d����DH���&�Zo�yvZ�z!l�/������)�Ķ<��N��?1(՚�!ļ��Y^H��bc��{q
N��ꍭ�@r3�<��{��-��7�K7�<V�Ϣ�v�{�
�1�L8G���r �'�O2��l�>��vhCy0�G�=�6@8q�aڤлkDF���^x~S0�����2�Ra$��ɑ��j~�\��	�����-��M>�֐j{|	�n�O��x��^ⅰ�n������O\ы��{�����ɭ�L-�&R��sm'�|�5f���!fc{�r`�����b�5_�L�=�4Yu/�CF��!�6�4y�������^,������a�&r��be�?� �2�n��}�#�D�3j��{	5h}QooL7qA�����ɧFQ�g<�gLW�S�to�"X&>))<hۇ琷B3�c6Mg!=�
V5߻�zb��D3X�1%�w�$��t}c��S�.3=G�|,IjG+�sS�l��B9�0��9��8;�K����-�k��5H�.��yV����\��"W��i$.]�[l?!�ao�y��#6?�6?;dF�fe�L���g��� >/>_���c�`��0�t>@:s��B��Y Li�;�n�l.3)I>��?_[�A��Y�Mq��?p0K|3�m��3=:��s}��9���.�źt "q6$��W";����o�5�YD��mSW�r����\�%�K�$��M	���b���!.ס.+1F�V�O�4��B��u�z�ڐ~y9�_NmxZ�oj��Aߪ�RW�Y��l�X�^����7V�|�3I�C��v��ٴ�Sg�8.;��\�MS����-��J�n�������IW�`
D�����d!QY)�0 ���r�A�k��*Vɟo�*�^ѓ��y��1bq�Ԝ�xLq��յ�����3M�$�l�Y�l-����d��:��c=��tq���n�`N�,���������b���M �4JyKb��O�}�"��5�j��~���:����,i>e�pL����5S�*��T�Obo�4-�^Ɋnk\���Ȕ
/ʩ7���p�w���5�����4>v�I>OX�Ƞ!���D��.'Գ����4oNm���V����Y���j�������
�Ŗ?���4s1~�&lyۚ��{*D+��C�Hڠ{�k׶Q�z�f`�f�����&�Q/��M��6����f�P��XPd�e1)�5�I�CZ�����:X�$�=l?�Xh��T���� ������?�ˀ�m���o����m}wP���
/���V�76S��Ó%7ʻ�b8�b�
`
M�;bP��b~S���C���9Iq�S- �>!�ƻ�e�>�'Q���Ӻ���]g�ᡑ<�جe@�AB"I�V���4�ҥ���w��eZ������ T���@�hEh}5��#�F���)m���L���Rf�iǌfJC�q�L{�yM���փ�8}K�zG��\fhͭ	#{����)yMo��Sl춭i'h�k��/9_D�XT|L����`��s�͡���^f�l�z��������N0��l�����j�o�9��Ξ��v���ӂ���T��%$�=�х����]��æ�c�eܻP�Y���ʼ���e�ꀣ��P��&��Ɍ��b[(]��|�[��(�4į���x��T��0�w�ixsLD.��HQ	��7��z�v4����s<s���gV���q��i�@�.w݄rX4�۲J��x����c�y.�u,O������jd�_�=r�ǅm�����+���7l_{������� �H�	N��+��O���L�K�(D:q�I\�~#�m�|���].��A�԰�H��sU����Ӭ.��x�Ի&V��|�t\>���	�t�l/�����L�І�湡� �����KU�S`��d�vb��Κ=�m��X{pp�㿘�\���cLv��R";H�d�2mJCݢ[��/���e�@�r����&S\>z)#^�sf5�eK��xb��@�ye��	���&[Bu�*&�%=�R�k����A{)5֏	&��8����[Y?��J�6�d$n�ǶQ�z��������f��8����6�K|taZ��t|J��rokG�#TT�3a��<�Uk���h�F�N'/T��@ɶ#���{��!'$\H� ��<VB"Ee���=�bM<�f�Z��>��7����;�6�K�zT3#c��[�;���d��Es|7�O���}�iն�9��P��@z\q��q�3����B�#���R��*v%S#�I�1+e׀w�&d~��P����*��eO��9��'Ť�|U:����4�g\s��n�b�H�|�ۼ�����ެ���SF�^���7�]4Q��S��t�k#� xa�t}�xH��jY�P��7���F���\��󋌝ڨ�5}"��7�@�h>l���W��{������rϐ���,={+ATQ;�w�;D�ŕ6� s��"R��8��̯�����gų�o]���d�P���N4EۥMc}��Mzmm�/ck'd��z[��_��>��� �� ��>�=��{[<W~̼sҐe�X/F�uq)������c9(��1�v�~ݢb��U���3�$��t��>��)N?h��v2o�B�?�~��>=3��uXi<t\?\�C���׷J2�V�01�Ȝ�Y9���w�K����~����t��~�=|�w�[n�{��MЃU����ig�JWU3�m-��Qʫ�Dp�z���&k�ޗ�ɯ}^�$ׁ^�@:���/`I�J{k��U��5�Rz�삧�$7X��B�U ��8ű�Y �]���~V�w�~L��w����a@:�G��m���CU=�f��s��+�;�-F�D:��=ň���[E�*�?����$�����IM`1��P���F�B%/�(LpA�o�t z�3Oެ5�G�����Ǆ��/I�~9�vꐽ�gWOd�� R�\5���'��8+�`f�ͤ� n��1E�BD�e}��_���;�>d����v�^��B��!�G����4��5�&�s���,��"u<��x3�ߑ����b~9n���>�.��%����#�T�\A�SV���.3����AYƤ�s�G(�����Fɭ�V�}�l���fCyM\��p�$ZÀ��d�?���=�֠�y��=���([�
|\-�E9�A& ����-�Z��ᨉ1��"`�쌟 b��TP^�qb0�<����C�F� ���j�P<���D���j�@��(������1z5shi:���|[�"/�\!���Fr�n�e�&Ǌ����!��у���C��G�`Yi�Y	(8����Ţ{�*dT�k�@05{%'���yX9�I��kggAu��צ�X:��F����	�?
mu6Ȫ��szy[m�����切�!r��2����K��S����奕�_P-��%YQ'k��/�Qsg0�nv�d%�%��)a�WU��#z��}r+̀��$?���P��s���R�r4 e	�H:yq��*���GJH�8@��l�oHᄩn�ێ9!}�n�����Ȃ2�d�	Q��h���;MB�'4���`ԼWIi ��8����2��oGʌe��g+��hw�Ut�8^�x���+�'���d����#�i�"�¾��FK6��z���Hw"콷H����r��K�J�X��q�R�yj����b/X@~����l�%PiiCp��r{ΆL:'c�hmtg(ϟZ�i`����+��iV�wX�z�������?���4�\�W����'$�T����RAral�ô3�xzj%P��J��hl钁K�@�]���~ ���L�I�J)��N��o{0qb�M� ��j���Ij�����m�jG�o/w�Y ���?KӒArϐ
d7�==����T�m&��X���f�eƆֿ��i�e�tV�%��Κq�C��}��p�1����F��0�X�}���l��)Q`͠�[j,������D�L����G#D#�J�垃k�+��T��2�d�J)�������GW]C��C7�TXHի��A�Rm,���i�lH���nbk�|��.D+�݋X�,����tч��X���X�Y>����I[Cfh��ƒuv�@�b��Z��a#����o	K���8-��{=���BIGe��`�[5��z-�o;�OD�E�*a����tFߦ��C�����,7.�ѳ�^sX1G��D/����2N+�B`RR���c�Ǘ���Hu�|�rA,a����o10��nK�1�LHBݿ�~َ>�y��C��W�2���V|����@�m��Z���V�3�i9'0����0d�c^M<O6�Wun���u�)Gҙ��,�J6��u��MX'�<�@��lQ��׮%\ӝ����X�jSi�5�$��0�\�Rr3+�$��U����t�xd���X�k���x6���_��f�����P�d�T8�����
)ߠ��T���h�L�P`	�U�h��#����R�	�r�۪���`�P��,!'V�:&(u�?<�TO�[��7�8��?j����!)��Im[)�I�J��Őg��N��qu�S��j���uL���F�I0
��`�K.�ʱ��;�m`�v|z��7�^�|Q�pyO�:���d{~�����(��I�뮮X�r����#yup�ɒgO^��̯�l|�>��t�Hk�^1Q��
$!Qʕ4i{��;�����(=(��w�]�.��u0�Qj|5��V�KiA;�T>��V�
J_�RSW�.����B� ��0�ፖT���Ė��޻�U�����/G���iήn����P0����9��K��01a?�ń����H�vJ7_��bP�B~U B�O6�V&L$Tg%0D�+&��?������@��\�0T ΃�}���F�N���W��$GpZ�xo�s
^gd M1��D���X��S@��o���djg�Oz�(���4�A�Y�������F)Sҍ��|0��:�Fk3�qjn�����9X*�Z�+�	�ZI'��V��ۂ���8D�������	�2��4��ͧV{�k����V��O9"����en���_6&� D��j4�tƥ�1kj�������3�T(�ֈ8��#��]�(�ܠ�D@���Um���������ŕ_T�\���P�v����o4����9�pJH���a�+NB���N%x�yr7,�V���1�o�Q�Λu��x���3Cs����#��-�~n����!qW/���&5�N�T�r�m&���&z�M�fe�z�4&di&k �c��Ƴu���}��|�������>�L�[:l �}JZ���s�.z�&w�8�%͞����BW��y>���[��m�
��%p���m�,[�(��)n�}ǂu�t�����cb�b�YFI�����K�X�)�Ȇ7�$��sх��?��O�ml'x�s��Q�,�!�MP�!�DU!�2�pN�>�2�����r�cheH嬔���,/�~�/k(^�:��'���p����P?�Eo���O�-t��]u����E�iw8`X��S����1� l?P.Ԋ��,�.�>QM�o��Z�x�Idr�#y`	Z�פ�ȏ� �^�o1��Sd��
x�2݅��i�!�?3h��.&��G�Ma�{{��_�Z�'����C+�1��:Dc�W�?u�C��K���x���b=5��ߎ�ݫR���5����.%��W��q������͂�f�o��;�b�)@T9��=_)�Q�y�ߝ��H����5����5�%12�'��l�|k>�����K�S�\�pv\�=�hw`J�A�&s�C�r�=��b p&�YF�zܿՈY�#�I�$δ�L
k�f�Uh�$9M��a޺��9_�����l�[�B��E��v���	�vaV՚6�#�]`�f�/�|�8�H�?�U#�.m�3|F�ny[K�ޭ��9�.��,��Lq	�g� ���������c�e(Il�`|�;�z���Q��k���=z2<BF�8`��Z7�-�.I�EŮ�QVI�ukK:�fϙ�!��i�t��gO:L57h�Q�;g޴Y&X�@41�����u|��N���ċ#�P1~k���x���jz&>�E- �?v�%o��r�#0Y�	d]+�m�v���z2�I�{��s�{��z�zG'X��<~Ǒ��w�S�Cugk��d�����c7�I_��8����������2��3��v>���dpg��+H'��K��L���VF~�������B^i4����ޡ�--��p;wW��5�sU���'٩H�೴�!^�O�WR\vQ����-p�P$¿���3��?@ &�G�!l�\'#f[����8�`L�@37Mc�=A>a��3]�������֗3R4�An��+�0g��%�	�j{��74�98|����Sq-%�JlQ��r��B�龰��/J^<�iX��3qP�^��1�un�e�@j2�Q������/����v�V�u}j�DYP�&��kDjzz���;|�7��jة�%d���'��\��bv�W�&�wp��i��s��p��e$� *�w+�@4�nլ��i��H6����V[��`=\f����5���vV+�k~�:3?/v\E�^�mR�	<qqOg�f��w���x�䐷���f�~�M��N�g�()QDE�U�����*��>2���!k&��Hi_�^s5ɣ��)N��#����l�Оj����Kns[s�r���m��&�+�/��D0��t�~;�Ϙ�p�َ�䀷�#�0Yg�3j�"�R�����-��:�Q���E9F�ױ���?12�Ts��"&�b"�1�b��θ�֊��b
¿��bF����\����@�#h�EoO�0���-�����{��n�r[߰!��]�`��Ef��jb�hC0�+�[�ߴ�VA+y���OkW��V֨�ڞ�`,�n?>��<�@�a�3�fof_��R;QB�>h���͒w���\�%��S�²�{��'h�$Z������s��� ���YvUC��7gѹ��"X�6�C���E[Q�B�d��c�u2P>�'��!�f'A��.sǬ��C���`�V.��`h�,������.� E���=�z��R��2�R���贊�>x��fվ؇���N�R��q��2����_�2B����x��tf��`xK��a��-$r*0��NK������� c�1^�{˯+Pf���u� >����j`E�Hϻ�E�%�;A�ֳsC[Wku�eGf�p]�愦�g�[�ږ|�r����/LQ�"c���8<�[s�X����̚AT���6)���pp|��Z��`���*g�e��߶t�}=���Q�����C�I����U�V%�h�j(������]�#��(����Re����YI����|5v����fAň^��N��,��H2����;�c��c�F݋���GɈ5T��A���Ͱ��&P�@�sn�?4�-�P�ԅO�*��Ƿ�֮�����PzEҶio�̟�w@�x�l$��� sv����D@�㵳���s)�D���G�͋���j[%j�&%�у�B�*0���`&�J�
���Q�������5]f1����/Z�
G��M�.-���(9V6I��;�z��O4��W��Ƥ���e��ј *1=!b�?���G����-��NC/�H�XS9C3�}��ɦJ䋓��Nu�r}� q�#_ 	˕e��GN�u��a(@|b4/)�����G��$t���8��%-��4�/��