��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���ohǫ�R�q͉L9��!Cj��!�_!,�ٔ�P�%���5^'�H������p�ϼ'/d�9�)���E��(܃�[�"�d7�+��Nm.a}����/�W�2��Cz]Њ2���X��w��t��P�{0櫢���d�B��{�B���*��M�L!�W�q��U�[��W���"M^x()
�$�v�����W�cu�Ic@���*E�z`�:8��Ҩ�׊�ݱ�ZU`��J����J�����Oۋ��ߤ�K_,�Ib����N�uU׵1{��S~.���z=yA�=��W�Bp�}�̋��%�_S\����Zՠ�,�fd�����Ul����҂�AC���71�Q�[Cs���$��@�骋�c�9�0���O��T8߅e����5�G����\����X�����kq��]4�P��c��q����0G�����(�x�x�bu ���տ����J�h�GBt��x�,)Zb�
��c�!޾bGI�� Q4+{[��P��&����AC}M\����&�����i�j��5�_�g��ރDt�:�o�P/$K]W�߇2kbQS�����Z�G����������]0)�7\���������.�K3���L����Pv]6�y���M�S̚�1�-�GVHT��~��pw�՟�,>�,�:nmn�	��VY=^�pꖏ�g�ӈ5v)��ڊ��Y�uu&���`�&8���t�\݁�73L�FGj�-�����l�� ����)?�߹�Q>��bn3��z�[���2W��U�����e��qv^�g�FDLG�a����-���f���b�����y����U�&:R%Ҧ����J�� lp<��U�Ϳ��ԃy�7�v2�x�ߖI�������G\�{�[D������搨��^Rt�<\7�s����2��E�*N_�eu�KZ�ƣ_d�F���w���
$O�]��Z�l�/�g84���T[�5���͏��1��p	.�ir�}f�@�C~U5�X� �J�݈3��`2z��k��Z���,ڱ�5:>@����/vh�.c6H#��7]��Z<,!��G㩪�)1�(�T�T���������>����V�GL����^ʤZ�۬/���b��̂���|5��-0�la��1>?*����1UQV���Y]�h2��U�Qې(��~���{�	���P?yۘ�W�Ä(Lh0�~���8ÐG������㎚�w�*���j$ fA�����RQ�f��g͓�:�KƯt�C�9姐�xgwJ�=��~�y��̂:��T*��e���6E�����}���OagS;h}�v6��zr9���G͋*kx/��f��f�� �+
X2��<���.Og��w3��N�^��D�
���)/�<����)z^g`��M`:�0���笣�f]=F]
M��ǵu���F�����Շ,-9C���\p-l�A5|7u�ر���Eg�uAE�8 VL�	e}
���e9[�\�R���cOV�ܙ����^e�4z�����I��;we����n���NG���8��ȇ���;<yh�waQ<B��E��~�������:*u���+�/B9��M��y�3a��ǸE�+!����Hr�4��B��&nrcژ2̡�X��+�\"���>�2��J��!r�H5����y�޺� 8{4��@e�D���E�$u�~��hn>˹�:.���<,��8�� :���j�{��i�TO�<��,

:���w��JX�R��x��%NoF�d?��9�?i|�f
�W�ɑ_  �JE³pL�����-�WQ�g��p��=ҩ>�f_����_Q�+��;L��z�!c�[|iC��U�8��4�~s&���n��޸& 2��J���Z�J���p��{��q2��h:�
):ޭP�c��(�������ÿ�;���%���E _��od֥�KM��.*��Z�GB
�|l�JW�	HL��4濤��ao�2uC枼��C\�����;̙�"ܣK�#�G��l�!_��8L��Ż��A�s�'�o��5��h�C^wͺ��n��͇�(	oI���&���7.�3��0���Q����m�9��H�`;�L��君�yhL�5�J�sD�L4D�b�	��5RC��>M���$�vCO�hH�z�߻��1�����<�,l�D��P��wq3�k\����?P�ʉ�;����v;sh|+\J�f�*�7d�6I:I �܋iN��<�]�ϓY���?sh$n�W_<Q@�.K~D�%�22����o@��i9ѥ"�{����Y�Q �O,0���QV�]��,�T':��oo8�l���(�(���n��6&��B+�^���Ɨ�Э������:M۫?���{`�Il�������0�Jj~�7�R�e��g�����*��	��hlJk���R)�W����`{�,����7����L�s�&�+)�]�ܯ�:���C�D��c���$�WZ_N�3B嵴�� 4p���k.��8�
�V����d�L�OX���0�����P	�(Fo�]�\�sjS�E��5�b�\/���?�2�i8�(�W�W
�d��� ��ejm6��� OE�#���	W���P�!��y�9�I1R�4�w$�7�X�Hq��>`|]��=6O妁���@��O��L�=���������P�oN��ϵ�|��ڸ��0yZHA�����o���u�����ċ�V�3�CV7*)o�����3;@C�A0a�\�ʨZ��e�l�c��q�̶��A�� 8�A�����x4�,/s7������(l���q��3[ː9�Y��B�g��+�2~b�~)��&1Pۻ$����u�~�=�[��|D�Z	�h�aqb⧲�@]��R������?�I/�3��q�Μ-��Ϛ�@fq�v�˴��}Y�np��b���l�)N�1�6�]��(���bd׼�ۉ���
�bS�-ئ��;c����㰅���P�p�����Bx�� �����Ai�7/7Y�Ե���^��˛%m�ŇZQ{-�O���F���'�o4��)�����,��[��c+L��\�v��E���o)a�/���E��~�"ԉ^���^,���e<�f֤��t��I��/qNG�������%�P�*��3���ˬ��X'��kEm<r����t�m�V^'8{f�b'v�I��^�c)�K�1v4����I�,,��+��3X�!L5�.5��InϮ��u��#��F�6�\���16rf~��>��F�-�Ï$������>�A��=�7�h�v4��7>���48O�%O�K� ��0�`1�[�!@�\�v��*�@l��S#zyҒ�����R}W�U�\4ͦ� X�HxL�%�z�ӷ��p�,a�gL��y�"��WJXڴ�W���P4W���ڪ���qnR�+��I���R�������.tŹg�SZ��&98n{��<��S�X�B���a�qs�����<�]��&�
�<�����5�L������AMC���$�!#s��C�qo�90Ѽc�����b�jU����(�d��[����l��:y)A�^l_�6��3�6�#mR��˾k\-����䄠�%Z�X	2,�-��m=+��%��^��
=p���6��yl�����%�T��#.��Q�x|�9�"�ȓ���� �;-wg�P�	F�L_��)�v�je��T��Β2~�v��#�2x��mX������M�STg��i��.L.���ֵ3c?τcԚ��yw1zDi����򗾪�0;��������Ӥ%�Eh�����,O@�s�����W��Wǯw1k2���Mp]���B��Q��KƦ���J%fR�1��+����}(�Yb�����y����l�k�8��	N���ek�>N��ByZZiU@�>��s)�e�b�(ũd�\����8!{%��P���?��լ+�ӊ�Dy����dk���+S��$�vU��N䓪n��n�N�1M�J|`z]:�̓O��a�W�4d�C��-�hm(ϼ'�#3�9,��0ɹx�a!|]&$��w=��+���Lv�+�@�i�~A�2�
�w���g� ��,:�)�=کq�#�;�7]����Ƭ.�^�����19��[���}��`���G��R�?������I'?E)K(
"]ۻ�^���릊ԵѪ�Q٤�G7LjD��)R_TI�|�y���ʀ��Q����گ�F�ک)4� �!3�t�`�%�L>��Y��?��&��R���@�+�b�,�7��eR��y���@$vP�	uqh�Z�+C��<h�I�\��y{��"�-���%V%9��DKw{@��L�Yd�[�׶)c�
,R� B��}��?w�P���T�\)�̞�L�7A� �r��R�e����A����~�:��_UN6J��n�*I��T��To"f��׶�6┨'*�n~E����w%~�|��
�Y����i+f~uM���꽩��N����Բ���=���&2y߽3sc����W{�h�E,)�i���d3.�����]U���U~4F*~�&��^��wx�h����9���Ɨ��=N���R+�R���|:�S'i���ڵ��.,ۏ�o����yfEb����D�ૣ	�T�����@3���#�~���2�1�U���C��k$z�e�I�x��t!D<#}b�h���ƶ�j��T�o�Y��b|K�4��αP#>����yW�g�M�:���>��%�ҧ�`FyX����/���A��O�(�.�� l�ۂV7]����$��x��p�]O�d�x�^�p��.�-�TX��͚��I�oˢya��̰��h�/���Vnow�Ve�Y�t�bb\��'B�3��J���s`�z�֣�	���I�o�ߕ�6�t��p�"Y�F�n�N��w
�RU����	5��|L�}��&�\
R��kI2%0�]��{�ɖ������u�s1{sm���ׄ���j���s$��`.X'�C�lq����KO?��ּ4�
�����W,�W��N9鯓N���1�-N>�-n�c���?p�A�0���,+S��p�E*��h�a-��L�Ӻ-��籧|���Po���2�A��$�����}�(�F�`7<�<�G�Z;������������;�]�4�!Gv}�1$��t�̚ ����Q��^�G�;���Os͌A'_���*wZ����r�S�d����`����MP�xҨ�9w���-n����چ �YS�_<v4���x"%G����/G��Bi��,�q��L~y����ќ%���x�'��9�!L^�:.ہ戮�x���R�uw}Gu�(g���+��:��lD^.��32��֒���V@��І��d��Y?�m�cYݺ�.�7����m�ª�����g"�J������E�v��d�~M�\3/��i��l����
�%�vj1�z{nw�fT�{uH��qg��-`��&��������>8{��'{��	��ZC,E�>�`5���J�7v��h��|<h�<,����E7�_b���.�/�½�	�ۉϪ:+oϝT�؝�ƭ-�����1��e<2�a��8��$z��ޠB�
ߑl�h���pUg�vO\��c�!��c�?� ѶQ|&Yb��ȗ��NH����R�wFkP"�K�*9�S��*�h��N�M�mL����o�ᨯ�ƱJ�JA������0LA*��JP�Ҙ
�:�5D�� 4����&��J-]w��F��cX�����#�6Nn����g���ߥ�@�~�$�m�͡9�a�O �B�����ASe9-+ҙ�B�+����<7������9��y������/Z�
���-cn�������[wZc����]��GB�M��K&���lu�8��k��o��H����m�vQN��:P����I
�GV��� ��nK���!Q)��j�$��a���uBjLY��ZͿE�≁c�� ��;i�w�Ǣ�!,;ئ�M�v�����Y~,���[�Ci��2�T��L�N/�U%
�u.p�@k�V���U�索I�`�@{����R����?�e�d!<���#��{�vE��N�_O��q0CE��&�K[��B�t	��7t�n�4��G;K'Y�|I%�$�3>�a0��*&`Ob!_��?Mr��3����hR���N�U׿�h��栨Ht���!$��A��:�qͳ+����CV���1�m7sCI7����҈�5C)3��֬F�f�ٞr�����3`�v�3�uI�s�9 �FUK��R�n�S�nE�R���O�����m��8�-��M��c���3��,��3�J�WIS���+�wGN�f�)V׭��C|#�ȑQ��(k��֊ə��^��z�����<��ɭ���O�>�[����Yq�l\J�������9�|�bgw��9� ��gw[��:�����)S. ��f�x�"B�D��}��w�:*	P�Rз�-�J�w�����B������-9g_q��{"~� �����&m�}�p)��D�u�����S��,��M�guq1F�`H,� 9��q�
o�,�-C�*Y����;"Ŵ�f�ef��D�	�3��)[��4�@����<���&�z*�n�oay�d�t��@�վ	�����se�y�
��B齨��u�3��%�o�%�V;���Lj�3WHg�{�?h��/t��Se�vF8�sk��8�;y�v%�����a�icQ߸p�|�(}ةa��5k��KK^t*��ͮ�L�`�狆8FG� ���@p��H_�<��Ȉ`�xXH�F��D��='�S�gUj���\J^��󲡹6+c`#�Q2�1��=����PJ6]���l|/P��*�r��*��ڹ2%��*�|�X��f�����>�˯ �?'℡ 9|Q`O�7��]���v������qET�yd�)6��$�ì���>g�
����C����+�ӭ�+z��?�-�S�H�"���T2Љvb�W�/�p�*
�|��;>�V�������P)k*|���e�
���NUn�
�cP�s߿D���vΔ��?hI&���X�����BÏ��cB|W����J���l������ؾ�C����0in&,}��A$��	K�O� /}����E�Ҍ���n7�
a�t\y�^���*�Е�
�Q�9�N��-�:�j�_
,�����+I�����d:�z��(�CNq��=���s�/5�n�?GFܓUt��4rӆ|*s�C�ͯ��s�o2 ��h��Ѵ���Ͽm���ۋ�I=FA�� l?L�ѭ���(|�BO eʖu�
����ģ���̡5ɰ�U���Z#Q#�' ����Ѷ��7�l���F�*K:�E/J�ua�+
�T���h���@�� Ą7��C��(��)t��s�Ws���!<�\�̙Մ
�5�[hleM��d�y�P햀�C.�3c1��f�`Q�b��v�� <�J�l^He�QK�
���ĴO��3?������jc/d5Yc����(�&�_T;�dQ\ѕ�3�=�q������?	�Jj:�OL�}m����b$2̾u�-HfL������4����aeJ���$i��/r�L��Ӿ���l��\���iu��O�������?��&c(߽<����6 �ƈ"�����ڮ6&>��a��h���M%�߃p��ڳ-,��BC�-����G��F��Z�F��s�,������7�MmzboX���1�m�@ʇ:�����=f��툪D���6#
�R7"|�+/�'F�Eql.��O#�*ܨ.�.�Q;��p(�)�Q�9�DbL����p<@�dÿ9�Z@?���_�u��;�A�Nt
TJ�0�c�e��a"�e���ĲN���	���}Oz����]`��N�7�U~��t��+{z;q>�Im�p+�ރ��M���Pe�@�O��2S�O��qݳr*o���ÇNʿ�
��3ײ�]�G11Hv� ��B�@�<���� �pHL�
vU��7�<ne0��ԮzNR�8�dx"�>C��+LK�\���s�^��>]�U�^P��'�
�W��r�`��,0��{�� /����7#X��5����=h�;H���H���s&'/�s�ݼ͡�9�l#�}��<��mm+��&b�qѳ�3�O�e��^�eC�[3m5����%,*Pae�F���K�<
�~c�& $����ntB�w���o|�S�nӹ!G��]����V�S0�l�x��V�/��/R7�3a�>��雎��z�͊k#95�6Ҳ�Â�n=�o�ǡ#J੓���2�@��Pٖ�N�]����Y|�q�;��ON�>a�t��.,�_>4,�%��v��`\���غb« �B=ޒd-X�r��ݻkR���ʐ��*HfH4'n�=%��d7�՘�c$�#��c�Ԙ1�&�1�������CJ`?�D����L*���������Xi|���zF�!9_���:7���ҨC6v�խ�U��v:��'���y���fPp]�[�dB(�������R5��G�S��������O7,��o6L��%�GA�3�	�T�(L`S��m�Q;?�Y6�SYK@�����Ԅ�9��K4�*�u�s���K}/�{c^H���z���w�i/}5O��4���Tj1i��h2��G98�%�(Cq�'��,76�n�A����d�В���x|�2P�|
r]�v $$�~�����e:ޮ�����d��7[�U��d8$"�[m�vt�fy�$� A�}��f�`$�j�9�xF��Ј6OV,���)GN�)%ɷ[�}�3�k��F���y�����=jD���7j`V���I��D��^R��4�~�iӑ�� 8�0M��O�)Ўf~�W����?��`܇G�v�7N��Z!g���v�ߝR,�f��7?��	z:m3����^�/����K&���:}�k�����E����#��pE��� �ᕁ;�Ûe�T�D��c!
d�-� S�8`���]��2�8���@�Ҏu jէ�?���u
�dKUFr;ې�`t�s`Ԉ`4����"f����.��~���z��sam�^���Ӡ�	�#�?���樓ӖSp��&����օ���d"-P�����x��'܉963���:�rt��B��S���[�lJ��^��6G�s�kM/�)��W��1�Վ��A�	U'�z�$�v�E�mi��C��B�~L6G�b�4&�kI�-����
��_��eMI�[����>.vVo����}����+�ec�=�������������e��B���ϯ�,x���ֶt�H�y^O��;��*��e�\"~=����5 !>������'9�G[�I�����u�6��XFFOTΔ�mh8-�qbpW���`�p8���P+ΰV��"3=�q�/ԟ��Z�k�9�W�1��:j��JY�z�� ï��F�`���X�}K̮x)6�3����A_�`����>%|�C#�cK��s�&���Ԯ#@�t�z,H�v=m��8�=u�L�A�p�R��ߗ|��Iۄܜ�F�隌]�e$�`��|pzi���V0�q�q��GO�����:[|��6����K�₁�F>�ŕʄ���ȻSCl7:����/X��fms�������o�w��ݝp,��X����l Ҏ"Ʋ���C��k����rs�	�j��;�&���W�B~#�f��ck���� �����hΧ���s���Xm�j�x�M)v��vy!3��_l
�=F�U}����.>B*�<>���I�����.��h	x[��a
����6#��;GS���I���BF�f���B�]�v�R4#��Z���b�HQ7��K���+���'ځ``!�E�D� ��y6�4Y���s�ݽ򑖛�� 
��@8"?��ం��P��ؔ�1�U�/��&��X��1xz���-���v��Z8�q��G.��9�.�N��d|F4�Nn'4����a��8�WK1�Y�Yg����|!DZI ��(#;�܆��i�p�)��<\S֬�8����`h�	�c�o�&hF�Q=��"��pUa�Yp*�P\n5��l�`��G�9kpM��lyF��'f�������)I���;{_���V�2��[���^d�=4��##rP�rB�~,��}Q*��<}���irn�+ίZ{�s�i�n���[|���~$�6fz^�X]��a��K��+�P�z�����Z��d2�\=�ވ��WmPG�~��1�ʫ�g���k'H�?*�P�]
#��pL��qv�R�_`��-�#W�^1�dEo��0K�PT�:h�j���\�{�T����7���vy!��fD�窙����O����b:��M��1��鴮�.��ʶdJ��GN��l�d��p4F�8�����s,t�7��x�4T�Yr�1@s�	<�#����Oy�Ժ�/�
N5��s �>�&ӏ�-��5��h�9Mr;�Ǒ�B��}i�w���i�cd�D1t@�F9vb���x�#i,���/�
Uw.vez4���%��'�&��2d�y����j�?�)fN��#�u�Ó���Kq��w1��u�@��<��zx��\�G}[4Gt�@���ș��	�r��jA{��P�	[~��Z_ƴ=�m�Y�i7c������5-
b�Fdly|xN���=�C�PW����t�A�@�"�_��Mt�~�9�x.�����$��y�3##k��)�ȫ�y�������xg\U����r<�!k���;q|B^l� h�`O��s`c���8�:K̈́�jD�+3R��l1ڄ�}D���kC�	HY���,����4�8X.��QH�	PfXcU�Dud������kS6���$.CW�z����hG�B�w:#����<-�E���9�\y�AI�\ ��Р���m���[��d��ĻZA����&O�T� bt�τ�{뎠4"2]��:�h_��?*�&6a���_�
4Y�Ȧ��O���[.�rd�4]��,y��x�ܒf��7� ��ϛ��JаL+jk���r��ZP�^Ǣ��x	���È��`�Z��;N�T��+���%i���\���D��նJ ���aY�rI�q=.�1Qb	��B�ˇ�(ĉ�92��X��鵬���]�IQ��w�\>x�zN�I�Ф`��L|ؤ�ø`Q���NF5�L�/p�����ڻ,���;�B�gӱYy�%��@(%&$�N[ �y^c��夲%�I�33YkvBS�F�x�y���c�Q�D�K�o$T!�/��� w��ם����c��#�2}m�@ޢ���a�ٓҩ:hcD���v�>}��{��{w2Ku7��^���n��=
��0cT���<�ӂ�~���-��Q����r���P�U��Nb�1*�� t��X�j�һ��Pfa�69�[�G�|6�g��l�����ۼ�0F]B�.��A����T��m��uqL�#]%�d��I'�=O���D*U��ʖ�`O<XEGf��ܪ-ƈ�;W�!22$�N��v�"��I�ޱI��3V�?]"� $�8����̶oC��|1 5l��6�ر����K|_�C=�R��F.����&�N	cᥥ��X��
��l�}�Ⱥ���yT7!���ՏP�PS����k奰�F�&@����cu�^;���'_�{F�,���G����`�J���n�T�w��-�083�iZP����<N#Z���F���Fهu���΂��2�roF�Ƽ������.�Ϯe�ݧ�U�>�$��|�l
�<oW���IN�'T��Z�4��qSc^<���$Y�93D�R�F�8�'�]#�h��w?enE����I(��B�x'!YK�V�<pR��]qۗ�x��eG=elD�SP+�W�j9Fj��@h��4κ�<O��ߚ�%���T�V���z���ti^��~�ӕ���{�Q��#�OU��8c�^Im(t�`A��v���U)�(���9��o�0����F-�Ai"x^l��cʆѾ.r�Nn��=��0\E�,`�7�� ���DM����S�fR�8��$j�⣐\�|(��ݓ%�g�wO���+\0i�f�"�k���agu�;��#x��@�o��wp������~0S>�$m@�_"�,�X���l������]_� %�8]�F�����1�w�!|�"�`V��M"vd�wdh3��ۊ�Vn}N@'�����q�lV����{�\�J�k¸ +��]^��;(h:�FQ4�g/l/)��a�"������Ueլ��"�/{�'��,x E�%����(n�&-F��W!P���(���0AW�t�0�v*r�������(���h��wJ*b���e�]l�����b9uZ�ٸJ!��{vP۰ H�w���q��h~W�J�[C��q�Q%ø¢zϠ���	t�
k���w����CV'�Qc���yw�Βyx��OI��)�P��w�Kz>�N���:��5{����	������tQCԶ�М���W���]N�s�w�uS]�>�͒�pM_�)<[��j���Nbϳ� P?g���/ANƧs��]L ;���R���8aAk2�"3l/�n̎ʤ$cje-�(���ҿ��K��7�T�e��&y�G�	n�9�������s�o�����^�۶�
;� ��f�T�7����I��\>��al�ϕ��'�ª��P�6�������#ъ��m@G�Q���OKĸe�a<&���� ��6��?�NI"�q %�|3fX� t��/uʑH)%�tD�:����m�+��M��!�G����:N�Gb���)�L`J"HWc���R��C�:���[ٷyv܂\
S��	�J,ZL���^Z��6��@�V��z_R��y��͔Q��^��E�-�1)0�Nf����7htp�'�R�(�V�[%�T�F�zqZ=��zr�Ԝn(u��|�fz���8����f���B�n��`�!\�~��c�|aټ��?��1u�!v��h�7"�wa���S*�q��#  ����!D���π;�K��a��Y���-�! ���R�NM8�]j���n(А��@D ���ݑi�*jC��H��D=V�`�uslY�R�hC-������X&�c$�P؀1� �t���MҐ]����+�T:�E���
�f�*��4�����#@0�ÕT���Ej�]�>{����zžI���M< �a�o��;���2|�33���Uόᏼ,e��u���T~@c��Y�ݦʉ�=�-������K<��u�
���PNP.��*�� �c#�ڏ�����)�#���g�i#�b�����A��&�c=&<]���k��Ш�㺦�hٚ*wt�!�>/����TO8�%�; �<F�t��Y�}kdg�j!��-�0�~�M"���h�=8N�ҡ��h�)q`B̒c�����3"���&���(���Gwگ2t�q�h��PW���Ҙ��f��rx��A	#�xǰ�\�X����)��AR�=OR�wy���^t',��vBsy���L��	P8���x+Ԟ�X����<,��_��i��e��(�8�QmL�-q$/�p;�26X�a�Y6ߡ
_*����SɆo��ɬ�![�u%�2	���O���yY��	��P��+D,�DU�Gt~-F�,	�n��4r. -ۓŁX�v��꺙�S���'��Kh��Z�tg���y�-�>�y�-�e�����s���/���õ�#{ژ�]r4�T�K���eڼ5�x���@gv�Ң%����K,�$mD7>u��3^����oG!�T��@��BO�$�jU>L��f�a �#��B���h1��;~�߆Ⱦ�N�֒�7=�U���WW�� �-'jL��tN]F�8o.X���S��Z�����XDZV�Y��?�6����zi'N�����ҭg�ɱE�1���s5������2d���A��H��u�4�>�\�Q�8�@Ӆ�|��'��9C׫���1>۾�e���[�Zf�Ew�I<<>��VڅN��ܹ.\^.f�R�I�.6�ZdZ5���QH�糤�����R��7�"�_��/�q/^Y����H�Az��(p[�"��9M�f�}��	%��M�lIM�p9��+B��`�)i���Ӽ��
onb(��Y|z��3༁o�T� ��?��u�B����q6�L`�� S�F$/��FV�Q3bl��^�$���Ç�ch^�֪V��s8� ��02�_S���p+{W~�U�	���v�ќRm�5���Q��g��ɧ#�<1�"�Wh�dd����ҏ�~c��!B�D��@�5��_�_,_�_�?��i�D��g�C�®�$sl�<�E/7���T(Yhn0��?�p����Co�w; ��M���J�w�\J�fS hZ��TgCqS�2O���c�[~
�?��O+X��!w�̟����<i�����=*�]&����"�0���C�70�6�����ϊƍC�=ILA����[�h=S}�D�:ĕ*qgm�.LΩXQ�WϚ����\f&�,|ڤW#����9<�. /mdᲕw���},2����nf2�lٔQ?;Y������q�{15�k��si�,7@t���i>�'MAQ^�?5�J�ɻ����aBi�X<��{�^��
;����4Ӟ�X�� :�ڴ�/2�.�cr\��UCZ�8��.#f�o8��l��	y�V�=υN���lrq���MeLW�-��(�kYA� �H@��nO��r�`��j��y��U6v�gE�|�G
<�G���@��sy��ɽ�hL`.��"*�A
	���wX�	<�G\�0)��;o\7%PjM�z�T�c���k��	��EhY�����4y�wjZu/��KO�"��j�C~WMV�z&4w[5��V��-�h����������nh�����7yow�-�y�2�+��Pz_\��K��`A�]vO��U�70`����ܻȘ��҂�%U�Y0�ؽ����ࢸqa3�9+B��nu~�]F <��p�>��N�o�x��"���m���ٔ�^S��?�/����U�%��rP�������05M�3"��/Rw�/��	��Iy��S���n�m���E��9�p��
I����10����O�����=��`j'|�[L06��m��Z��(�dy��X���s}��<��m� ���4�@\�A>�J��ir=���6��J�zJ����T.�����r�z�=&���"����~���0��(��-.z����T����q���Nm>�iR�	|4$����0���㨂�Rk���ےa�f? �#>q0q[ ݩ�B �;]���y����b<0��/�E;_4�1 �=Z�����O䰄=D	�Яd*QI��ۓB����m��hZ���gʅ!9l>�Q)g�t�,����[���Ė���i�{��H�W�	l}'4�خ���uNI��B�\6Ck��e�þ����j܌_�E�z�-���t�)���p�3?Ǫ�5f�k�_R9�x�eŎQ?�~?��w��r���o�������`d�Pe�h�A??��eY��D��흖�e��'�a[%v`'O�$�l��u&�y�EL��J�hY���-<�p�z�ÔB]i˞t,�1IP��T��.���K1K&��ceG�����ב�8�D �h��z�,�qr�U�v�[�$t��`��B��[h�:Xc:���|32d��a3k��(��#�}��"�_�і�=�f��{\6������9X�R��S�3�w�^*�oT).�JC`�y�0�<oc�=�[���(�����ko��$��{���B��{�[d���FJ�p���Һ�B�[��}�?�����V�!�[Pʭ�,��S��¼��dU|��U@`�������U�����¯�c�ҭ��l�K>����֤��ZX��%Z<M�0ƪeA�3(���ɪ�F���o���M3�ٯ��mSX�/�)��"� `΍�"���>b��45LkW)R�yG���TB?�)�'����*�y�_���n�W�_CL�`~����&�}����+���A�f�ᨡ��~^�ݼ��rQ�1�9�1Q�;y�P�㫗��dq��"�O>�u[5���I\��>a�\1Z8��s�2�|��J���C8�l���{V`�Ʈ��@���a�I��G�D���K�Ɂ.�5�4rj��&
��`�~N��DrlՆ��q�����)����k4��~��I
��)I�
��["sr��eo�zxJwR�Y�h���7[-6�|�у���������~�kZΕ^�)U^"j:|�%���enG�}o�{jW����gO6s:�ŬZ9<������ CM��0G,��z�9�ێWu�L�Y��mf�kr��)��P��b����%��i|8}�U��w	�7����k�f� ��?��ki��TC�U�p'��	v�Jϰ߄O��F�vg��)��	 tR|�k�޾��V�12�v�kP�Bէ�Ur�t����(��$����*�ڶ4M���BRO�Ǡ�4+'�=���a�3c��=;�ef2��7��$O�P�#D��M���y8�,�P���h��?�J� �c�lDT^*�|	5
}�#����0�	b*�F�\xQ֗�"��-bv���Xe�,r�1|�s��)A����
R���֬��~4�%P�B��K��m�{�=���Xa���v�1�S";�^���ṌyYb{H¡�Ofn[���s̓���iO�, ��A�ynЀ�r�B�a
 &X���z�«�a��l?�%�P<��؄OKz���c��&�d/aF�d�/īK��&`ߠyh?�H�4�x^�XG]U��t�}
dh��3��m��TΝo���.6i'��(ܩ>����l\��9�7��r�L����8s+�rl�e�߫��9�N��"��+���[��ӆ�x����;_�+C�~�� 돋(��)
(����d��y������y�o�x����L�Ic���n8a�8�f��r�V��%��3iѷE�˒B<9Y@�L���	A��p�y-���Q���w�|��Ü��,8�
�\A�P�Sl���J&G��;ǤG�"�A�QU�My���ӄ��A1Y��z>�H�Ky-wkn��G9���~��g�9��a�'SW����}df�3Ci�텸�Vފ��6K.'����q8��e��� ��%����('`(�}G���8zF[����������{`��w9�ߵI�o�ƪ